-- soc_system.vhd

-- Generated using ACDS version 20.1 711

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity soc_system is
	port (
		ad1939_abclk_clk                    : in    std_logic                     := '0';             --            ad1939_abclk.clk
		ad1939_alrclk_clk                   : in    std_logic                     := '0';             --           ad1939_alrclk.clk
		ad1939_mclk_clk                     : in    std_logic                     := '0';             --             ad1939_mclk.clk
		ad1939_physical_asdata2             : in    std_logic                     := '0';             --         ad1939_physical.asdata2
		ad1939_physical_dbclk               : out   std_logic;                                        --                        .dbclk
		ad1939_physical_dlrclk              : out   std_logic;                                        --                        .dlrclk
		ad1939_physical_dsdata1             : out   std_logic;                                        --                        .dsdata1
		clk_clk                             : in    std_logic                     := '0';             --                     clk.clk
		hps_f2h_cold_reset_req_reset_n      : in    std_logic                     := '0';             --  hps_f2h_cold_reset_req.reset_n
		hps_f2h_debug_reset_req_reset_n     : in    std_logic                     := '0';             -- hps_f2h_debug_reset_req.reset_n
		hps_f2h_warm_reset_req_reset_n      : in    std_logic                     := '0';             --  hps_f2h_warm_reset_req.reset_n
		hps_h2f_reset_reset_n               : out   std_logic;                                        --           hps_h2f_reset.reset_n
		hps_hps_io_hps_io_emac1_inst_TX_CLK : out   std_logic;                                        --              hps_hps_io.hps_io_emac1_inst_TX_CLK
		hps_hps_io_hps_io_emac1_inst_TXD0   : out   std_logic;                                        --                        .hps_io_emac1_inst_TXD0
		hps_hps_io_hps_io_emac1_inst_TXD1   : out   std_logic;                                        --                        .hps_io_emac1_inst_TXD1
		hps_hps_io_hps_io_emac1_inst_TXD2   : out   std_logic;                                        --                        .hps_io_emac1_inst_TXD2
		hps_hps_io_hps_io_emac1_inst_TXD3   : out   std_logic;                                        --                        .hps_io_emac1_inst_TXD3
		hps_hps_io_hps_io_emac1_inst_RXD0   : in    std_logic                     := '0';             --                        .hps_io_emac1_inst_RXD0
		hps_hps_io_hps_io_emac1_inst_MDIO   : inout std_logic                     := '0';             --                        .hps_io_emac1_inst_MDIO
		hps_hps_io_hps_io_emac1_inst_MDC    : out   std_logic;                                        --                        .hps_io_emac1_inst_MDC
		hps_hps_io_hps_io_emac1_inst_RX_CTL : in    std_logic                     := '0';             --                        .hps_io_emac1_inst_RX_CTL
		hps_hps_io_hps_io_emac1_inst_TX_CTL : out   std_logic;                                        --                        .hps_io_emac1_inst_TX_CTL
		hps_hps_io_hps_io_emac1_inst_RX_CLK : in    std_logic                     := '0';             --                        .hps_io_emac1_inst_RX_CLK
		hps_hps_io_hps_io_emac1_inst_RXD1   : in    std_logic                     := '0';             --                        .hps_io_emac1_inst_RXD1
		hps_hps_io_hps_io_emac1_inst_RXD2   : in    std_logic                     := '0';             --                        .hps_io_emac1_inst_RXD2
		hps_hps_io_hps_io_emac1_inst_RXD3   : in    std_logic                     := '0';             --                        .hps_io_emac1_inst_RXD3
		hps_hps_io_hps_io_sdio_inst_CMD     : inout std_logic                     := '0';             --                        .hps_io_sdio_inst_CMD
		hps_hps_io_hps_io_sdio_inst_D0      : inout std_logic                     := '0';             --                        .hps_io_sdio_inst_D0
		hps_hps_io_hps_io_sdio_inst_D1      : inout std_logic                     := '0';             --                        .hps_io_sdio_inst_D1
		hps_hps_io_hps_io_sdio_inst_CLK     : out   std_logic;                                        --                        .hps_io_sdio_inst_CLK
		hps_hps_io_hps_io_sdio_inst_D2      : inout std_logic                     := '0';             --                        .hps_io_sdio_inst_D2
		hps_hps_io_hps_io_sdio_inst_D3      : inout std_logic                     := '0';             --                        .hps_io_sdio_inst_D3
		hps_hps_io_hps_io_usb1_inst_D0      : inout std_logic                     := '0';             --                        .hps_io_usb1_inst_D0
		hps_hps_io_hps_io_usb1_inst_D1      : inout std_logic                     := '0';             --                        .hps_io_usb1_inst_D1
		hps_hps_io_hps_io_usb1_inst_D2      : inout std_logic                     := '0';             --                        .hps_io_usb1_inst_D2
		hps_hps_io_hps_io_usb1_inst_D3      : inout std_logic                     := '0';             --                        .hps_io_usb1_inst_D3
		hps_hps_io_hps_io_usb1_inst_D4      : inout std_logic                     := '0';             --                        .hps_io_usb1_inst_D4
		hps_hps_io_hps_io_usb1_inst_D5      : inout std_logic                     := '0';             --                        .hps_io_usb1_inst_D5
		hps_hps_io_hps_io_usb1_inst_D6      : inout std_logic                     := '0';             --                        .hps_io_usb1_inst_D6
		hps_hps_io_hps_io_usb1_inst_D7      : inout std_logic                     := '0';             --                        .hps_io_usb1_inst_D7
		hps_hps_io_hps_io_usb1_inst_CLK     : in    std_logic                     := '0';             --                        .hps_io_usb1_inst_CLK
		hps_hps_io_hps_io_usb1_inst_STP     : out   std_logic;                                        --                        .hps_io_usb1_inst_STP
		hps_hps_io_hps_io_usb1_inst_DIR     : in    std_logic                     := '0';             --                        .hps_io_usb1_inst_DIR
		hps_hps_io_hps_io_usb1_inst_NXT     : in    std_logic                     := '0';             --                        .hps_io_usb1_inst_NXT
		hps_hps_io_hps_io_spim1_inst_CLK    : out   std_logic;                                        --                        .hps_io_spim1_inst_CLK
		hps_hps_io_hps_io_spim1_inst_MOSI   : out   std_logic;                                        --                        .hps_io_spim1_inst_MOSI
		hps_hps_io_hps_io_spim1_inst_MISO   : in    std_logic                     := '0';             --                        .hps_io_spim1_inst_MISO
		hps_hps_io_hps_io_spim1_inst_SS0    : out   std_logic;                                        --                        .hps_io_spim1_inst_SS0
		hps_hps_io_hps_io_uart0_inst_RX     : in    std_logic                     := '0';             --                        .hps_io_uart0_inst_RX
		hps_hps_io_hps_io_uart0_inst_TX     : out   std_logic;                                        --                        .hps_io_uart0_inst_TX
		hps_hps_io_hps_io_i2c1_inst_SDA     : inout std_logic                     := '0';             --                        .hps_io_i2c1_inst_SDA
		hps_hps_io_hps_io_i2c1_inst_SCL     : inout std_logic                     := '0';             --                        .hps_io_i2c1_inst_SCL
		hps_hps_io_hps_io_gpio_inst_GPIO09  : inout std_logic                     := '0';             --                        .hps_io_gpio_inst_GPIO09
		hps_hps_io_hps_io_gpio_inst_GPIO35  : inout std_logic                     := '0';             --                        .hps_io_gpio_inst_GPIO35
		hps_hps_io_hps_io_gpio_inst_GPIO40  : inout std_logic                     := '0';             --                        .hps_io_gpio_inst_GPIO40
		hps_hps_io_hps_io_gpio_inst_GPIO53  : inout std_logic                     := '0';             --                        .hps_io_gpio_inst_GPIO53
		hps_hps_io_hps_io_gpio_inst_GPIO54  : inout std_logic                     := '0';             --                        .hps_io_gpio_inst_GPIO54
		hps_hps_io_hps_io_gpio_inst_GPIO61  : inout std_logic                     := '0';             --                        .hps_io_gpio_inst_GPIO61
		hps_i2c0_out_data                   : out   std_logic;                                        --                hps_i2c0.out_data
		hps_i2c0_sda                        : in    std_logic                     := '0';             --                        .sda
		hps_i2c0_clk_clk                    : out   std_logic;                                        --            hps_i2c0_clk.clk
		hps_i2c0_scl_in_clk                 : in    std_logic                     := '0';             --         hps_i2c0_scl_in.clk
		hps_spim0_txd                       : out   std_logic;                                        --               hps_spim0.txd
		hps_spim0_rxd                       : in    std_logic                     := '0';             --                        .rxd
		hps_spim0_ss_in_n                   : in    std_logic                     := '0';             --                        .ss_in_n
		hps_spim0_ssi_oe_n                  : out   std_logic;                                        --                        .ssi_oe_n
		hps_spim0_ss_0_n                    : out   std_logic;                                        --                        .ss_0_n
		hps_spim0_ss_1_n                    : out   std_logic;                                        --                        .ss_1_n
		hps_spim0_ss_2_n                    : out   std_logic;                                        --                        .ss_2_n
		hps_spim0_ss_3_n                    : out   std_logic;                                        --                        .ss_3_n
		hps_spim0_sclk_out_clk              : out   std_logic;                                        --      hps_spim0_sclk_out.clk
		memory_mem_a                        : out   std_logic_vector(14 downto 0);                    --                  memory.mem_a
		memory_mem_ba                       : out   std_logic_vector(2 downto 0);                     --                        .mem_ba
		memory_mem_ck                       : out   std_logic;                                        --                        .mem_ck
		memory_mem_ck_n                     : out   std_logic;                                        --                        .mem_ck_n
		memory_mem_cke                      : out   std_logic;                                        --                        .mem_cke
		memory_mem_cs_n                     : out   std_logic;                                        --                        .mem_cs_n
		memory_mem_ras_n                    : out   std_logic;                                        --                        .mem_ras_n
		memory_mem_cas_n                    : out   std_logic;                                        --                        .mem_cas_n
		memory_mem_we_n                     : out   std_logic;                                        --                        .mem_we_n
		memory_mem_reset_n                  : out   std_logic;                                        --                        .mem_reset_n
		memory_mem_dq                       : inout std_logic_vector(31 downto 0) := (others => '0'); --                        .mem_dq
		memory_mem_dqs                      : inout std_logic_vector(3 downto 0)  := (others => '0'); --                        .mem_dqs
		memory_mem_dqs_n                    : inout std_logic_vector(3 downto 0)  := (others => '0'); --                        .mem_dqs_n
		memory_mem_odt                      : out   std_logic;                                        --                        .mem_odt
		memory_mem_dm                       : out   std_logic_vector(3 downto 0);                     --                        .mem_dm
		memory_oct_rzqin                    : in    std_logic                     := '0';             --                        .oct_rzqin
		reset_reset_n                       : in    std_logic                     := '0'              --                   reset.reset_n
	);
end entity soc_system;

architecture rtl of soc_system is
	component AD1939_hps_audio_mini is
		port (
			sys_clk            : in  std_logic                     := 'X';             -- clk
			sys_reset          : in  std_logic                     := 'X';             -- reset
			AD1939_ADC_ABCLK   : in  std_logic                     := 'X';             -- clk
			AD1939_ADC_ALRCLK  : in  std_logic                     := 'X';             -- clk
			AD1939_ADC_channel : out std_logic_vector(1 downto 0);                     -- channel
			AD1939_ADC_data    : out std_logic_vector(31 downto 0);                    -- data
			AD1939_ADC_error   : out std_logic_vector(1 downto 0);                     -- error
			AD1939_ADC_valid   : out std_logic;                                        -- valid
			AD1939_DAC_channel : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- channel
			AD1939_DAC_data    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- data
			AD1939_DAC_error   : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- error
			AD1939_DAC_valid   : in  std_logic                     := 'X';             -- valid
			AD1939_ADC_ASDATA2 : in  std_logic                     := 'X';             -- asdata2
			AD1939_DAC_DBCLK   : out std_logic;                                        -- dbclk
			AD1939_DAC_DLRCLK  : out std_logic;                                        -- dlrclk
			AD1939_DAC_DSDATA1 : out std_logic                                         -- dsdata1
		);
	end component AD1939_hps_audio_mini;

	component soc_system_PLL_using_AD1939_MCLK is
		port (
			refclk   : in  std_logic := 'X'; -- clk
			rst      : in  std_logic := 'X'; -- reset
			outclk_0 : out std_logic;        -- clk
			locked   : out std_logic         -- export
		);
	end component soc_system_PLL_using_AD1939_MCLK;

	component soc_system_SystemID is
		port (
			clock    : in  std_logic                     := 'X'; -- clk
			reset_n  : in  std_logic                     := 'X'; -- reset_n
			readdata : out std_logic_vector(31 downto 0);        -- readdata
			address  : in  std_logic                     := 'X'  -- address
		);
	end component soc_system_SystemID;

	component soc_system_hps is
		generic (
			F2S_Width : integer := 2;
			S2F_Width : integer := 2
		);
		port (
			h2f_cold_rst_n           : out   std_logic;                                         -- reset_n
			f2h_cold_rst_req_n       : in    std_logic                      := 'X';             -- reset_n
			f2h_dbg_rst_req_n        : in    std_logic                      := 'X';             -- reset_n
			f2h_warm_rst_req_n       : in    std_logic                      := 'X';             -- reset_n
			spim0_txd                : out   std_logic;                                         -- txd
			spim0_rxd                : in    std_logic                      := 'X';             -- rxd
			spim0_ss_in_n            : in    std_logic                      := 'X';             -- ss_in_n
			spim0_ssi_oe_n           : out   std_logic;                                         -- ssi_oe_n
			spim0_ss_0_n             : out   std_logic;                                         -- ss_0_n
			spim0_ss_1_n             : out   std_logic;                                         -- ss_1_n
			spim0_ss_2_n             : out   std_logic;                                         -- ss_2_n
			spim0_ss_3_n             : out   std_logic;                                         -- ss_3_n
			spim0_sclk_out           : out   std_logic;                                         -- clk
			i2c0_scl                 : in    std_logic                      := 'X';             -- clk
			i2c0_out_clk             : out   std_logic;                                         -- clk
			i2c0_out_data            : out   std_logic;                                         -- out_data
			i2c0_sda                 : in    std_logic                      := 'X';             -- sda
			mem_a                    : out   std_logic_vector(14 downto 0);                     -- mem_a
			mem_ba                   : out   std_logic_vector(2 downto 0);                      -- mem_ba
			mem_ck                   : out   std_logic;                                         -- mem_ck
			mem_ck_n                 : out   std_logic;                                         -- mem_ck_n
			mem_cke                  : out   std_logic;                                         -- mem_cke
			mem_cs_n                 : out   std_logic;                                         -- mem_cs_n
			mem_ras_n                : out   std_logic;                                         -- mem_ras_n
			mem_cas_n                : out   std_logic;                                         -- mem_cas_n
			mem_we_n                 : out   std_logic;                                         -- mem_we_n
			mem_reset_n              : out   std_logic;                                         -- mem_reset_n
			mem_dq                   : inout std_logic_vector(31 downto 0)  := (others => 'X'); -- mem_dq
			mem_dqs                  : inout std_logic_vector(3 downto 0)   := (others => 'X'); -- mem_dqs
			mem_dqs_n                : inout std_logic_vector(3 downto 0)   := (others => 'X'); -- mem_dqs_n
			mem_odt                  : out   std_logic;                                         -- mem_odt
			mem_dm                   : out   std_logic_vector(3 downto 0);                      -- mem_dm
			oct_rzqin                : in    std_logic                      := 'X';             -- oct_rzqin
			hps_io_emac1_inst_TX_CLK : out   std_logic;                                         -- hps_io_emac1_inst_TX_CLK
			hps_io_emac1_inst_TXD0   : out   std_logic;                                         -- hps_io_emac1_inst_TXD0
			hps_io_emac1_inst_TXD1   : out   std_logic;                                         -- hps_io_emac1_inst_TXD1
			hps_io_emac1_inst_TXD2   : out   std_logic;                                         -- hps_io_emac1_inst_TXD2
			hps_io_emac1_inst_TXD3   : out   std_logic;                                         -- hps_io_emac1_inst_TXD3
			hps_io_emac1_inst_RXD0   : in    std_logic                      := 'X';             -- hps_io_emac1_inst_RXD0
			hps_io_emac1_inst_MDIO   : inout std_logic                      := 'X';             -- hps_io_emac1_inst_MDIO
			hps_io_emac1_inst_MDC    : out   std_logic;                                         -- hps_io_emac1_inst_MDC
			hps_io_emac1_inst_RX_CTL : in    std_logic                      := 'X';             -- hps_io_emac1_inst_RX_CTL
			hps_io_emac1_inst_TX_CTL : out   std_logic;                                         -- hps_io_emac1_inst_TX_CTL
			hps_io_emac1_inst_RX_CLK : in    std_logic                      := 'X';             -- hps_io_emac1_inst_RX_CLK
			hps_io_emac1_inst_RXD1   : in    std_logic                      := 'X';             -- hps_io_emac1_inst_RXD1
			hps_io_emac1_inst_RXD2   : in    std_logic                      := 'X';             -- hps_io_emac1_inst_RXD2
			hps_io_emac1_inst_RXD3   : in    std_logic                      := 'X';             -- hps_io_emac1_inst_RXD3
			hps_io_sdio_inst_CMD     : inout std_logic                      := 'X';             -- hps_io_sdio_inst_CMD
			hps_io_sdio_inst_D0      : inout std_logic                      := 'X';             -- hps_io_sdio_inst_D0
			hps_io_sdio_inst_D1      : inout std_logic                      := 'X';             -- hps_io_sdio_inst_D1
			hps_io_sdio_inst_CLK     : out   std_logic;                                         -- hps_io_sdio_inst_CLK
			hps_io_sdio_inst_D2      : inout std_logic                      := 'X';             -- hps_io_sdio_inst_D2
			hps_io_sdio_inst_D3      : inout std_logic                      := 'X';             -- hps_io_sdio_inst_D3
			hps_io_usb1_inst_D0      : inout std_logic                      := 'X';             -- hps_io_usb1_inst_D0
			hps_io_usb1_inst_D1      : inout std_logic                      := 'X';             -- hps_io_usb1_inst_D1
			hps_io_usb1_inst_D2      : inout std_logic                      := 'X';             -- hps_io_usb1_inst_D2
			hps_io_usb1_inst_D3      : inout std_logic                      := 'X';             -- hps_io_usb1_inst_D3
			hps_io_usb1_inst_D4      : inout std_logic                      := 'X';             -- hps_io_usb1_inst_D4
			hps_io_usb1_inst_D5      : inout std_logic                      := 'X';             -- hps_io_usb1_inst_D5
			hps_io_usb1_inst_D6      : inout std_logic                      := 'X';             -- hps_io_usb1_inst_D6
			hps_io_usb1_inst_D7      : inout std_logic                      := 'X';             -- hps_io_usb1_inst_D7
			hps_io_usb1_inst_CLK     : in    std_logic                      := 'X';             -- hps_io_usb1_inst_CLK
			hps_io_usb1_inst_STP     : out   std_logic;                                         -- hps_io_usb1_inst_STP
			hps_io_usb1_inst_DIR     : in    std_logic                      := 'X';             -- hps_io_usb1_inst_DIR
			hps_io_usb1_inst_NXT     : in    std_logic                      := 'X';             -- hps_io_usb1_inst_NXT
			hps_io_spim1_inst_CLK    : out   std_logic;                                         -- hps_io_spim1_inst_CLK
			hps_io_spim1_inst_MOSI   : out   std_logic;                                         -- hps_io_spim1_inst_MOSI
			hps_io_spim1_inst_MISO   : in    std_logic                      := 'X';             -- hps_io_spim1_inst_MISO
			hps_io_spim1_inst_SS0    : out   std_logic;                                         -- hps_io_spim1_inst_SS0
			hps_io_uart0_inst_RX     : in    std_logic                      := 'X';             -- hps_io_uart0_inst_RX
			hps_io_uart0_inst_TX     : out   std_logic;                                         -- hps_io_uart0_inst_TX
			hps_io_i2c1_inst_SDA     : inout std_logic                      := 'X';             -- hps_io_i2c1_inst_SDA
			hps_io_i2c1_inst_SCL     : inout std_logic                      := 'X';             -- hps_io_i2c1_inst_SCL
			hps_io_gpio_inst_GPIO09  : inout std_logic                      := 'X';             -- hps_io_gpio_inst_GPIO09
			hps_io_gpio_inst_GPIO35  : inout std_logic                      := 'X';             -- hps_io_gpio_inst_GPIO35
			hps_io_gpio_inst_GPIO40  : inout std_logic                      := 'X';             -- hps_io_gpio_inst_GPIO40
			hps_io_gpio_inst_GPIO53  : inout std_logic                      := 'X';             -- hps_io_gpio_inst_GPIO53
			hps_io_gpio_inst_GPIO54  : inout std_logic                      := 'X';             -- hps_io_gpio_inst_GPIO54
			hps_io_gpio_inst_GPIO61  : inout std_logic                      := 'X';             -- hps_io_gpio_inst_GPIO61
			h2f_rst_n                : out   std_logic;                                         -- reset_n
			h2f_axi_clk              : in    std_logic                      := 'X';             -- clk
			h2f_AWID                 : out   std_logic_vector(11 downto 0);                     -- awid
			h2f_AWADDR               : out   std_logic_vector(29 downto 0);                     -- awaddr
			h2f_AWLEN                : out   std_logic_vector(3 downto 0);                      -- awlen
			h2f_AWSIZE               : out   std_logic_vector(2 downto 0);                      -- awsize
			h2f_AWBURST              : out   std_logic_vector(1 downto 0);                      -- awburst
			h2f_AWLOCK               : out   std_logic_vector(1 downto 0);                      -- awlock
			h2f_AWCACHE              : out   std_logic_vector(3 downto 0);                      -- awcache
			h2f_AWPROT               : out   std_logic_vector(2 downto 0);                      -- awprot
			h2f_AWVALID              : out   std_logic;                                         -- awvalid
			h2f_AWREADY              : in    std_logic                      := 'X';             -- awready
			h2f_WID                  : out   std_logic_vector(11 downto 0);                     -- wid
			h2f_WDATA                : out   std_logic_vector(63 downto 0);                     -- wdata
			h2f_WSTRB                : out   std_logic_vector(7 downto 0);                      -- wstrb
			h2f_WLAST                : out   std_logic;                                         -- wlast
			h2f_WVALID               : out   std_logic;                                         -- wvalid
			h2f_WREADY               : in    std_logic                      := 'X';             -- wready
			h2f_BID                  : in    std_logic_vector(11 downto 0)  := (others => 'X'); -- bid
			h2f_BRESP                : in    std_logic_vector(1 downto 0)   := (others => 'X'); -- bresp
			h2f_BVALID               : in    std_logic                      := 'X';             -- bvalid
			h2f_BREADY               : out   std_logic;                                         -- bready
			h2f_ARID                 : out   std_logic_vector(11 downto 0);                     -- arid
			h2f_ARADDR               : out   std_logic_vector(29 downto 0);                     -- araddr
			h2f_ARLEN                : out   std_logic_vector(3 downto 0);                      -- arlen
			h2f_ARSIZE               : out   std_logic_vector(2 downto 0);                      -- arsize
			h2f_ARBURST              : out   std_logic_vector(1 downto 0);                      -- arburst
			h2f_ARLOCK               : out   std_logic_vector(1 downto 0);                      -- arlock
			h2f_ARCACHE              : out   std_logic_vector(3 downto 0);                      -- arcache
			h2f_ARPROT               : out   std_logic_vector(2 downto 0);                      -- arprot
			h2f_ARVALID              : out   std_logic;                                         -- arvalid
			h2f_ARREADY              : in    std_logic                      := 'X';             -- arready
			h2f_RID                  : in    std_logic_vector(11 downto 0)  := (others => 'X'); -- rid
			h2f_RDATA                : in    std_logic_vector(63 downto 0)  := (others => 'X'); -- rdata
			h2f_RRESP                : in    std_logic_vector(1 downto 0)   := (others => 'X'); -- rresp
			h2f_RLAST                : in    std_logic                      := 'X';             -- rlast
			h2f_RVALID               : in    std_logic                      := 'X';             -- rvalid
			h2f_RREADY               : out   std_logic;                                         -- rready
			f2h_axi_clk              : in    std_logic                      := 'X';             -- clk
			f2h_AWID                 : in    std_logic_vector(7 downto 0)   := (others => 'X'); -- awid
			f2h_AWADDR               : in    std_logic_vector(31 downto 0)  := (others => 'X'); -- awaddr
			f2h_AWLEN                : in    std_logic_vector(3 downto 0)   := (others => 'X'); -- awlen
			f2h_AWSIZE               : in    std_logic_vector(2 downto 0)   := (others => 'X'); -- awsize
			f2h_AWBURST              : in    std_logic_vector(1 downto 0)   := (others => 'X'); -- awburst
			f2h_AWLOCK               : in    std_logic_vector(1 downto 0)   := (others => 'X'); -- awlock
			f2h_AWCACHE              : in    std_logic_vector(3 downto 0)   := (others => 'X'); -- awcache
			f2h_AWPROT               : in    std_logic_vector(2 downto 0)   := (others => 'X'); -- awprot
			f2h_AWVALID              : in    std_logic                      := 'X';             -- awvalid
			f2h_AWREADY              : out   std_logic;                                         -- awready
			f2h_AWUSER               : in    std_logic_vector(4 downto 0)   := (others => 'X'); -- awuser
			f2h_WID                  : in    std_logic_vector(7 downto 0)   := (others => 'X'); -- wid
			f2h_WDATA                : in    std_logic_vector(127 downto 0) := (others => 'X'); -- wdata
			f2h_WSTRB                : in    std_logic_vector(15 downto 0)  := (others => 'X'); -- wstrb
			f2h_WLAST                : in    std_logic                      := 'X';             -- wlast
			f2h_WVALID               : in    std_logic                      := 'X';             -- wvalid
			f2h_WREADY               : out   std_logic;                                         -- wready
			f2h_BID                  : out   std_logic_vector(7 downto 0);                      -- bid
			f2h_BRESP                : out   std_logic_vector(1 downto 0);                      -- bresp
			f2h_BVALID               : out   std_logic;                                         -- bvalid
			f2h_BREADY               : in    std_logic                      := 'X';             -- bready
			f2h_ARID                 : in    std_logic_vector(7 downto 0)   := (others => 'X'); -- arid
			f2h_ARADDR               : in    std_logic_vector(31 downto 0)  := (others => 'X'); -- araddr
			f2h_ARLEN                : in    std_logic_vector(3 downto 0)   := (others => 'X'); -- arlen
			f2h_ARSIZE               : in    std_logic_vector(2 downto 0)   := (others => 'X'); -- arsize
			f2h_ARBURST              : in    std_logic_vector(1 downto 0)   := (others => 'X'); -- arburst
			f2h_ARLOCK               : in    std_logic_vector(1 downto 0)   := (others => 'X'); -- arlock
			f2h_ARCACHE              : in    std_logic_vector(3 downto 0)   := (others => 'X'); -- arcache
			f2h_ARPROT               : in    std_logic_vector(2 downto 0)   := (others => 'X'); -- arprot
			f2h_ARVALID              : in    std_logic                      := 'X';             -- arvalid
			f2h_ARREADY              : out   std_logic;                                         -- arready
			f2h_ARUSER               : in    std_logic_vector(4 downto 0)   := (others => 'X'); -- aruser
			f2h_RID                  : out   std_logic_vector(7 downto 0);                      -- rid
			f2h_RDATA                : out   std_logic_vector(127 downto 0);                    -- rdata
			f2h_RRESP                : out   std_logic_vector(1 downto 0);                      -- rresp
			f2h_RLAST                : out   std_logic;                                         -- rlast
			f2h_RVALID               : out   std_logic;                                         -- rvalid
			f2h_RREADY               : in    std_logic                      := 'X';             -- rready
			h2f_lw_axi_clk           : in    std_logic                      := 'X';             -- clk
			h2f_lw_AWID              : out   std_logic_vector(11 downto 0);                     -- awid
			h2f_lw_AWADDR            : out   std_logic_vector(20 downto 0);                     -- awaddr
			h2f_lw_AWLEN             : out   std_logic_vector(3 downto 0);                      -- awlen
			h2f_lw_AWSIZE            : out   std_logic_vector(2 downto 0);                      -- awsize
			h2f_lw_AWBURST           : out   std_logic_vector(1 downto 0);                      -- awburst
			h2f_lw_AWLOCK            : out   std_logic_vector(1 downto 0);                      -- awlock
			h2f_lw_AWCACHE           : out   std_logic_vector(3 downto 0);                      -- awcache
			h2f_lw_AWPROT            : out   std_logic_vector(2 downto 0);                      -- awprot
			h2f_lw_AWVALID           : out   std_logic;                                         -- awvalid
			h2f_lw_AWREADY           : in    std_logic                      := 'X';             -- awready
			h2f_lw_WID               : out   std_logic_vector(11 downto 0);                     -- wid
			h2f_lw_WDATA             : out   std_logic_vector(31 downto 0);                     -- wdata
			h2f_lw_WSTRB             : out   std_logic_vector(3 downto 0);                      -- wstrb
			h2f_lw_WLAST             : out   std_logic;                                         -- wlast
			h2f_lw_WVALID            : out   std_logic;                                         -- wvalid
			h2f_lw_WREADY            : in    std_logic                      := 'X';             -- wready
			h2f_lw_BID               : in    std_logic_vector(11 downto 0)  := (others => 'X'); -- bid
			h2f_lw_BRESP             : in    std_logic_vector(1 downto 0)   := (others => 'X'); -- bresp
			h2f_lw_BVALID            : in    std_logic                      := 'X';             -- bvalid
			h2f_lw_BREADY            : out   std_logic;                                         -- bready
			h2f_lw_ARID              : out   std_logic_vector(11 downto 0);                     -- arid
			h2f_lw_ARADDR            : out   std_logic_vector(20 downto 0);                     -- araddr
			h2f_lw_ARLEN             : out   std_logic_vector(3 downto 0);                      -- arlen
			h2f_lw_ARSIZE            : out   std_logic_vector(2 downto 0);                      -- arsize
			h2f_lw_ARBURST           : out   std_logic_vector(1 downto 0);                      -- arburst
			h2f_lw_ARLOCK            : out   std_logic_vector(1 downto 0);                      -- arlock
			h2f_lw_ARCACHE           : out   std_logic_vector(3 downto 0);                      -- arcache
			h2f_lw_ARPROT            : out   std_logic_vector(2 downto 0);                      -- arprot
			h2f_lw_ARVALID           : out   std_logic;                                         -- arvalid
			h2f_lw_ARREADY           : in    std_logic                      := 'X';             -- arready
			h2f_lw_RID               : in    std_logic_vector(11 downto 0)  := (others => 'X'); -- rid
			h2f_lw_RDATA             : in    std_logic_vector(31 downto 0)  := (others => 'X'); -- rdata
			h2f_lw_RRESP             : in    std_logic_vector(1 downto 0)   := (others => 'X'); -- rresp
			h2f_lw_RLAST             : in    std_logic                      := 'X';             -- rlast
			h2f_lw_RVALID            : in    std_logic                      := 'X';             -- rvalid
			h2f_lw_RREADY            : out   std_logic;                                         -- rready
			f2h_irq_p0               : in    std_logic_vector(31 downto 0)  := (others => 'X'); -- irq
			f2h_irq_p1               : in    std_logic_vector(31 downto 0)  := (others => 'X')  -- irq
		);
	end component soc_system_hps;

	component soc_system_jtag_uart is
		port (
			clk            : in  std_logic                     := 'X';             -- clk
			rst_n          : in  std_logic                     := 'X';             -- reset_n
			av_chipselect  : in  std_logic                     := 'X';             -- chipselect
			av_address     : in  std_logic                     := 'X';             -- address
			av_read_n      : in  std_logic                     := 'X';             -- read_n
			av_readdata    : out std_logic_vector(31 downto 0);                    -- readdata
			av_write_n     : in  std_logic                     := 'X';             -- write_n
			av_writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			av_waitrequest : out std_logic;                                        -- waitrequest
			av_irq         : out std_logic                                         -- irq
		);
	end component soc_system_jtag_uart;

	component soc_system_master_0 is
		generic (
			USE_PLI     : integer := 0;
			PLI_PORT    : integer := 50000;
			FIFO_DEPTHS : integer := 2
		);
		port (
			clk_clk              : in  std_logic                     := 'X';             -- clk
			clk_reset_reset      : in  std_logic                     := 'X';             -- reset
			master_address       : out std_logic_vector(31 downto 0);                    -- address
			master_readdata      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			master_read          : out std_logic;                                        -- read
			master_write         : out std_logic;                                        -- write
			master_writedata     : out std_logic_vector(31 downto 0);                    -- writedata
			master_waitrequest   : in  std_logic                     := 'X';             -- waitrequest
			master_readdatavalid : in  std_logic                     := 'X';             -- readdatavalid
			master_byteenable    : out std_logic_vector(3 downto 0);                     -- byteenable
			master_reset_reset   : out std_logic                                         -- reset
		);
	end component soc_system_master_0;

	component soc_system_onchip_memory is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			address    : in  std_logic_vector(12 downto 0) := (others => 'X'); -- address
			clken      : in  std_logic                     := 'X';             -- clken
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write      : in  std_logic                     := 'X';             -- write
			readdata   : out std_logic_vector(63 downto 0);                    -- readdata
			writedata  : in  std_logic_vector(63 downto 0) := (others => 'X'); -- writedata
			byteenable : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- byteenable
			reset      : in  std_logic                     := 'X';             -- reset
			reset_req  : in  std_logic                     := 'X';             -- reset_req
			freeze     : in  std_logic                     := 'X'              -- freeze
		);
	end component soc_system_onchip_memory;

	component pFIR_Testing_dataplane_avalon is
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			avalon_sink_valid        : in  std_logic                     := 'X';             -- valid
			avalon_sink_data         : in  std_logic_vector(31 downto 0) := (others => 'X'); -- data
			avalon_sink_channel      : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- channel
			avalon_sink_error        : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- error
			avalon_source_valid      : out std_logic;                                        -- valid
			avalon_source_data       : out std_logic_vector(31 downto 0);                    -- data
			avalon_source_channel    : out std_logic_vector(1 downto 0);                     -- channel
			avalon_source_error      : out std_logic_vector(1 downto 0);                     -- error
			avalon_slave_0_address   : in  std_logic                     := 'X';             -- address
			avalon_slave_0_read      : in  std_logic                     := 'X';             -- read
			avalon_slave_0_readdata  : out std_logic_vector(31 downto 0);                    -- readdata
			avalon_slave_0_write     : in  std_logic                     := 'X';             -- write
			avalon_slave_0_writedata : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			avalon_slave_1_address   : in  std_logic_vector(8 downto 0)  := (others => 'X'); -- address
			avalon_slave_1_read      : in  std_logic                     := 'X';             -- read
			avalon_slave_1_readdata  : out std_logic_vector(31 downto 0);                    -- readdata
			avalon_slave_1_write     : in  std_logic                     := 'X';             -- write
			avalon_slave_1_writedata : in  std_logic_vector(31 downto 0) := (others => 'X')  -- writedata
		);
	end component pFIR_Testing_dataplane_avalon;

	component soc_system_mm_interconnect_0 is
		port (
			hps_h2f_axi_master_awid                                        : in  std_logic_vector(11 downto 0) := (others => 'X'); -- awid
			hps_h2f_axi_master_awaddr                                      : in  std_logic_vector(29 downto 0) := (others => 'X'); -- awaddr
			hps_h2f_axi_master_awlen                                       : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- awlen
			hps_h2f_axi_master_awsize                                      : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- awsize
			hps_h2f_axi_master_awburst                                     : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- awburst
			hps_h2f_axi_master_awlock                                      : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- awlock
			hps_h2f_axi_master_awcache                                     : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- awcache
			hps_h2f_axi_master_awprot                                      : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- awprot
			hps_h2f_axi_master_awvalid                                     : in  std_logic                     := 'X';             -- awvalid
			hps_h2f_axi_master_awready                                     : out std_logic;                                        -- awready
			hps_h2f_axi_master_wid                                         : in  std_logic_vector(11 downto 0) := (others => 'X'); -- wid
			hps_h2f_axi_master_wdata                                       : in  std_logic_vector(63 downto 0) := (others => 'X'); -- wdata
			hps_h2f_axi_master_wstrb                                       : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- wstrb
			hps_h2f_axi_master_wlast                                       : in  std_logic                     := 'X';             -- wlast
			hps_h2f_axi_master_wvalid                                      : in  std_logic                     := 'X';             -- wvalid
			hps_h2f_axi_master_wready                                      : out std_logic;                                        -- wready
			hps_h2f_axi_master_bid                                         : out std_logic_vector(11 downto 0);                    -- bid
			hps_h2f_axi_master_bresp                                       : out std_logic_vector(1 downto 0);                     -- bresp
			hps_h2f_axi_master_bvalid                                      : out std_logic;                                        -- bvalid
			hps_h2f_axi_master_bready                                      : in  std_logic                     := 'X';             -- bready
			hps_h2f_axi_master_arid                                        : in  std_logic_vector(11 downto 0) := (others => 'X'); -- arid
			hps_h2f_axi_master_araddr                                      : in  std_logic_vector(29 downto 0) := (others => 'X'); -- araddr
			hps_h2f_axi_master_arlen                                       : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- arlen
			hps_h2f_axi_master_arsize                                      : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- arsize
			hps_h2f_axi_master_arburst                                     : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- arburst
			hps_h2f_axi_master_arlock                                      : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- arlock
			hps_h2f_axi_master_arcache                                     : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- arcache
			hps_h2f_axi_master_arprot                                      : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- arprot
			hps_h2f_axi_master_arvalid                                     : in  std_logic                     := 'X';             -- arvalid
			hps_h2f_axi_master_arready                                     : out std_logic;                                        -- arready
			hps_h2f_axi_master_rid                                         : out std_logic_vector(11 downto 0);                    -- rid
			hps_h2f_axi_master_rdata                                       : out std_logic_vector(63 downto 0);                    -- rdata
			hps_h2f_axi_master_rresp                                       : out std_logic_vector(1 downto 0);                     -- rresp
			hps_h2f_axi_master_rlast                                       : out std_logic;                                        -- rlast
			hps_h2f_axi_master_rvalid                                      : out std_logic;                                        -- rvalid
			hps_h2f_axi_master_rready                                      : in  std_logic                     := 'X';             -- rready
			clk_hps_clk_clk                                                : in  std_logic                     := 'X';             -- clk
			hps_h2f_axi_master_agent_clk_reset_reset_bridge_in_reset_reset : in  std_logic                     := 'X';             -- reset
			onchip_memory_reset1_reset_bridge_in_reset_reset               : in  std_logic                     := 'X';             -- reset
			onchip_memory_s1_address                                       : out std_logic_vector(12 downto 0);                    -- address
			onchip_memory_s1_write                                         : out std_logic;                                        -- write
			onchip_memory_s1_readdata                                      : in  std_logic_vector(63 downto 0) := (others => 'X'); -- readdata
			onchip_memory_s1_writedata                                     : out std_logic_vector(63 downto 0);                    -- writedata
			onchip_memory_s1_byteenable                                    : out std_logic_vector(7 downto 0);                     -- byteenable
			onchip_memory_s1_chipselect                                    : out std_logic;                                        -- chipselect
			onchip_memory_s1_clken                                         : out std_logic                                         -- clken
		);
	end component soc_system_mm_interconnect_0;

	component soc_system_mm_interconnect_1 is
		port (
			hps_h2f_lw_axi_master_awid                                        : in  std_logic_vector(11 downto 0) := (others => 'X'); -- awid
			hps_h2f_lw_axi_master_awaddr                                      : in  std_logic_vector(20 downto 0) := (others => 'X'); -- awaddr
			hps_h2f_lw_axi_master_awlen                                       : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- awlen
			hps_h2f_lw_axi_master_awsize                                      : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- awsize
			hps_h2f_lw_axi_master_awburst                                     : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- awburst
			hps_h2f_lw_axi_master_awlock                                      : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- awlock
			hps_h2f_lw_axi_master_awcache                                     : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- awcache
			hps_h2f_lw_axi_master_awprot                                      : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- awprot
			hps_h2f_lw_axi_master_awvalid                                     : in  std_logic                     := 'X';             -- awvalid
			hps_h2f_lw_axi_master_awready                                     : out std_logic;                                        -- awready
			hps_h2f_lw_axi_master_wid                                         : in  std_logic_vector(11 downto 0) := (others => 'X'); -- wid
			hps_h2f_lw_axi_master_wdata                                       : in  std_logic_vector(31 downto 0) := (others => 'X'); -- wdata
			hps_h2f_lw_axi_master_wstrb                                       : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- wstrb
			hps_h2f_lw_axi_master_wlast                                       : in  std_logic                     := 'X';             -- wlast
			hps_h2f_lw_axi_master_wvalid                                      : in  std_logic                     := 'X';             -- wvalid
			hps_h2f_lw_axi_master_wready                                      : out std_logic;                                        -- wready
			hps_h2f_lw_axi_master_bid                                         : out std_logic_vector(11 downto 0);                    -- bid
			hps_h2f_lw_axi_master_bresp                                       : out std_logic_vector(1 downto 0);                     -- bresp
			hps_h2f_lw_axi_master_bvalid                                      : out std_logic;                                        -- bvalid
			hps_h2f_lw_axi_master_bready                                      : in  std_logic                     := 'X';             -- bready
			hps_h2f_lw_axi_master_arid                                        : in  std_logic_vector(11 downto 0) := (others => 'X'); -- arid
			hps_h2f_lw_axi_master_araddr                                      : in  std_logic_vector(20 downto 0) := (others => 'X'); -- araddr
			hps_h2f_lw_axi_master_arlen                                       : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- arlen
			hps_h2f_lw_axi_master_arsize                                      : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- arsize
			hps_h2f_lw_axi_master_arburst                                     : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- arburst
			hps_h2f_lw_axi_master_arlock                                      : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- arlock
			hps_h2f_lw_axi_master_arcache                                     : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- arcache
			hps_h2f_lw_axi_master_arprot                                      : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- arprot
			hps_h2f_lw_axi_master_arvalid                                     : in  std_logic                     := 'X';             -- arvalid
			hps_h2f_lw_axi_master_arready                                     : out std_logic;                                        -- arready
			hps_h2f_lw_axi_master_rid                                         : out std_logic_vector(11 downto 0);                    -- rid
			hps_h2f_lw_axi_master_rdata                                       : out std_logic_vector(31 downto 0);                    -- rdata
			hps_h2f_lw_axi_master_rresp                                       : out std_logic_vector(1 downto 0);                     -- rresp
			hps_h2f_lw_axi_master_rlast                                       : out std_logic;                                        -- rlast
			hps_h2f_lw_axi_master_rvalid                                      : out std_logic;                                        -- rvalid
			hps_h2f_lw_axi_master_rready                                      : in  std_logic                     := 'X';             -- rready
			clk_hps_clk_clk                                                   : in  std_logic                     := 'X';             -- clk
			PLL_using_AD1939_MCLK_outclk0_clk                                 : in  std_logic                     := 'X';             -- clk
			hps_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset_reset : in  std_logic                     := 'X';             -- reset
			jtag_uart_reset_reset_bridge_in_reset_reset                       : in  std_logic                     := 'X';             -- reset
			master_0_clk_reset_reset_bridge_in_reset_reset                    : in  std_logic                     := 'X';             -- reset
			pFIR_Testing_0_reset_reset_bridge_in_reset_reset                  : in  std_logic                     := 'X';             -- reset
			SystemID_reset_reset_bridge_in_reset_reset                        : in  std_logic                     := 'X';             -- reset
			master_0_master_address                                           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- address
			master_0_master_waitrequest                                       : out std_logic;                                        -- waitrequest
			master_0_master_byteenable                                        : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			master_0_master_read                                              : in  std_logic                     := 'X';             -- read
			master_0_master_readdata                                          : out std_logic_vector(31 downto 0);                    -- readdata
			master_0_master_readdatavalid                                     : out std_logic;                                        -- readdatavalid
			master_0_master_write                                             : in  std_logic                     := 'X';             -- write
			master_0_master_writedata                                         : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			jtag_uart_avalon_jtag_slave_address                               : out std_logic_vector(0 downto 0);                     -- address
			jtag_uart_avalon_jtag_slave_write                                 : out std_logic;                                        -- write
			jtag_uart_avalon_jtag_slave_read                                  : out std_logic;                                        -- read
			jtag_uart_avalon_jtag_slave_readdata                              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			jtag_uart_avalon_jtag_slave_writedata                             : out std_logic_vector(31 downto 0);                    -- writedata
			jtag_uart_avalon_jtag_slave_waitrequest                           : in  std_logic                     := 'X';             -- waitrequest
			jtag_uart_avalon_jtag_slave_chipselect                            : out std_logic;                                        -- chipselect
			pFIR_Testing_0_avalon_slave_0_address                             : out std_logic_vector(0 downto 0);                     -- address
			pFIR_Testing_0_avalon_slave_0_write                               : out std_logic;                                        -- write
			pFIR_Testing_0_avalon_slave_0_read                                : out std_logic;                                        -- read
			pFIR_Testing_0_avalon_slave_0_readdata                            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			pFIR_Testing_0_avalon_slave_0_writedata                           : out std_logic_vector(31 downto 0);                    -- writedata
			pFIR_Testing_0_avalon_slave_1_address                             : out std_logic_vector(8 downto 0);                     -- address
			pFIR_Testing_0_avalon_slave_1_write                               : out std_logic;                                        -- write
			pFIR_Testing_0_avalon_slave_1_read                                : out std_logic;                                        -- read
			pFIR_Testing_0_avalon_slave_1_readdata                            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			pFIR_Testing_0_avalon_slave_1_writedata                           : out std_logic_vector(31 downto 0);                    -- writedata
			SystemID_control_slave_address                                    : out std_logic_vector(0 downto 0);                     -- address
			SystemID_control_slave_readdata                                   : in  std_logic_vector(31 downto 0) := (others => 'X')  -- readdata
		);
	end component soc_system_mm_interconnect_1;

	component soc_system_irq_mapper is
		port (
			clk           : in  std_logic                     := 'X'; -- clk
			reset         : in  std_logic                     := 'X'; -- reset
			receiver0_irq : in  std_logic                     := 'X'; -- irq
			sender_irq    : out std_logic_vector(31 downto 0)         -- irq
		);
	end component soc_system_irq_mapper;

	component soc_system_irq_mapper_001 is
		port (
			clk        : in  std_logic                     := 'X'; -- clk
			reset      : in  std_logic                     := 'X'; -- reset
			sender_irq : out std_logic_vector(31 downto 0)         -- irq
		);
	end component soc_system_irq_mapper_001;

	component soc_system_avalon_st_adapter is
		generic (
			inBitsPerSymbol : integer := 8;
			inUsePackets    : integer := 0;
			inDataWidth     : integer := 8;
			inChannelWidth  : integer := 3;
			inErrorWidth    : integer := 2;
			inUseEmptyPort  : integer := 0;
			inUseValid      : integer := 1;
			inUseReady      : integer := 1;
			inReadyLatency  : integer := 0;
			outDataWidth    : integer := 32;
			outChannelWidth : integer := 3;
			outErrorWidth   : integer := 2;
			outUseEmptyPort : integer := 0;
			outUseValid     : integer := 1;
			outUseReady     : integer := 1;
			outReadyLatency : integer := 0
		);
		port (
			in_clk_0_clk   : in  std_logic                     := 'X';             -- clk
			in_rst_0_reset : in  std_logic                     := 'X';             -- reset
			in_0_data      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- data
			in_0_valid     : in  std_logic                     := 'X';             -- valid
			in_0_error     : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- error
			in_0_channel   : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- channel
			out_0_data     : out std_logic_vector(31 downto 0);                    -- data
			out_0_valid    : out std_logic;                                        -- valid
			out_0_error    : out std_logic_vector(1 downto 0);                     -- error
			out_0_channel  : out std_logic_vector(1 downto 0)                      -- channel
		);
	end component soc_system_avalon_st_adapter;

	component soc_system_avalon_st_adapter_001 is
		generic (
			inBitsPerSymbol : integer := 8;
			inUsePackets    : integer := 0;
			inDataWidth     : integer := 8;
			inChannelWidth  : integer := 3;
			inErrorWidth    : integer := 2;
			inUseEmptyPort  : integer := 0;
			inUseValid      : integer := 1;
			inUseReady      : integer := 1;
			inReadyLatency  : integer := 0;
			outDataWidth    : integer := 32;
			outChannelWidth : integer := 3;
			outErrorWidth   : integer := 2;
			outUseEmptyPort : integer := 0;
			outUseValid     : integer := 1;
			outUseReady     : integer := 1;
			outReadyLatency : integer := 0
		);
		port (
			in_clk_0_clk   : in  std_logic                     := 'X';             -- clk
			in_rst_0_reset : in  std_logic                     := 'X';             -- reset
			in_0_data      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- data
			in_0_valid     : in  std_logic                     := 'X';             -- valid
			in_0_error     : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- error
			in_0_channel   : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- channel
			out_0_data     : out std_logic_vector(31 downto 0);                    -- data
			out_0_valid    : out std_logic;                                        -- valid
			out_0_error    : out std_logic_vector(1 downto 0);                     -- error
			out_0_channel  : out std_logic_vector(1 downto 0)                      -- channel
		);
	end component soc_system_avalon_st_adapter_001;

	component soc_system_rst_controller is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset_in0.reset
			clk            : in  std_logic := 'X'; --       clk.clk
			reset_out      : out std_logic;        -- reset_out.reset
			reset_in1      : in  std_logic := 'X';
			reset_in10     : in  std_logic := 'X';
			reset_in11     : in  std_logic := 'X';
			reset_in12     : in  std_logic := 'X';
			reset_in13     : in  std_logic := 'X';
			reset_in14     : in  std_logic := 'X';
			reset_in15     : in  std_logic := 'X';
			reset_in2      : in  std_logic := 'X';
			reset_in3      : in  std_logic := 'X';
			reset_in4      : in  std_logic := 'X';
			reset_in5      : in  std_logic := 'X';
			reset_in6      : in  std_logic := 'X';
			reset_in7      : in  std_logic := 'X';
			reset_in8      : in  std_logic := 'X';
			reset_in9      : in  std_logic := 'X';
			reset_req      : out std_logic;
			reset_req_in0  : in  std_logic := 'X';
			reset_req_in1  : in  std_logic := 'X';
			reset_req_in10 : in  std_logic := 'X';
			reset_req_in11 : in  std_logic := 'X';
			reset_req_in12 : in  std_logic := 'X';
			reset_req_in13 : in  std_logic := 'X';
			reset_req_in14 : in  std_logic := 'X';
			reset_req_in15 : in  std_logic := 'X';
			reset_req_in2  : in  std_logic := 'X';
			reset_req_in3  : in  std_logic := 'X';
			reset_req_in4  : in  std_logic := 'X';
			reset_req_in5  : in  std_logic := 'X';
			reset_req_in6  : in  std_logic := 'X';
			reset_req_in7  : in  std_logic := 'X';
			reset_req_in8  : in  std_logic := 'X';
			reset_req_in9  : in  std_logic := 'X'
		);
	end component soc_system_rst_controller;

	component soc_system_rst_controller_001 is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset_in0.reset
			clk            : in  std_logic := 'X'; --       clk.clk
			reset_out      : out std_logic;        -- reset_out.reset
			reset_req      : out std_logic;        --          .reset_req
			reset_in1      : in  std_logic := 'X';
			reset_in10     : in  std_logic := 'X';
			reset_in11     : in  std_logic := 'X';
			reset_in12     : in  std_logic := 'X';
			reset_in13     : in  std_logic := 'X';
			reset_in14     : in  std_logic := 'X';
			reset_in15     : in  std_logic := 'X';
			reset_in2      : in  std_logic := 'X';
			reset_in3      : in  std_logic := 'X';
			reset_in4      : in  std_logic := 'X';
			reset_in5      : in  std_logic := 'X';
			reset_in6      : in  std_logic := 'X';
			reset_in7      : in  std_logic := 'X';
			reset_in8      : in  std_logic := 'X';
			reset_in9      : in  std_logic := 'X';
			reset_req_in0  : in  std_logic := 'X';
			reset_req_in1  : in  std_logic := 'X';
			reset_req_in10 : in  std_logic := 'X';
			reset_req_in11 : in  std_logic := 'X';
			reset_req_in12 : in  std_logic := 'X';
			reset_req_in13 : in  std_logic := 'X';
			reset_req_in14 : in  std_logic := 'X';
			reset_req_in15 : in  std_logic := 'X';
			reset_req_in2  : in  std_logic := 'X';
			reset_req_in3  : in  std_logic := 'X';
			reset_req_in4  : in  std_logic := 'X';
			reset_req_in5  : in  std_logic := 'X';
			reset_req_in6  : in  std_logic := 'X';
			reset_req_in7  : in  std_logic := 'X';
			reset_req_in8  : in  std_logic := 'X';
			reset_req_in9  : in  std_logic := 'X'
		);
	end component soc_system_rst_controller_001;

	component soc_system_rst_controller_002 is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset_in0.reset
			reset_in1      : in  std_logic := 'X'; -- reset_in1.reset
			clk            : in  std_logic := 'X'; --       clk.clk
			reset_out      : out std_logic;        -- reset_out.reset
			reset_in10     : in  std_logic := 'X';
			reset_in11     : in  std_logic := 'X';
			reset_in12     : in  std_logic := 'X';
			reset_in13     : in  std_logic := 'X';
			reset_in14     : in  std_logic := 'X';
			reset_in15     : in  std_logic := 'X';
			reset_in2      : in  std_logic := 'X';
			reset_in3      : in  std_logic := 'X';
			reset_in4      : in  std_logic := 'X';
			reset_in5      : in  std_logic := 'X';
			reset_in6      : in  std_logic := 'X';
			reset_in7      : in  std_logic := 'X';
			reset_in8      : in  std_logic := 'X';
			reset_in9      : in  std_logic := 'X';
			reset_req      : out std_logic;
			reset_req_in0  : in  std_logic := 'X';
			reset_req_in1  : in  std_logic := 'X';
			reset_req_in10 : in  std_logic := 'X';
			reset_req_in11 : in  std_logic := 'X';
			reset_req_in12 : in  std_logic := 'X';
			reset_req_in13 : in  std_logic := 'X';
			reset_req_in14 : in  std_logic := 'X';
			reset_req_in15 : in  std_logic := 'X';
			reset_req_in2  : in  std_logic := 'X';
			reset_req_in3  : in  std_logic := 'X';
			reset_req_in4  : in  std_logic := 'X';
			reset_req_in5  : in  std_logic := 'X';
			reset_req_in6  : in  std_logic := 'X';
			reset_req_in7  : in  std_logic := 'X';
			reset_req_in8  : in  std_logic := 'X';
			reset_req_in9  : in  std_logic := 'X'
		);
	end component soc_system_rst_controller_002;

	signal hps_h2f_reset_reset                                           : std_logic;                     -- hps:h2f_rst_n -> [hps_h2f_reset_reset_n, hps_h2f_reset_reset_n:in]
	signal pll_using_ad1939_mclk_outclk0_clk                             : std_logic;                     -- PLL_using_AD1939_MCLK:outclk_0 -> [FE_Qsys_AD1939_Audio_Mini_v1_0:sys_clk, avalon_st_adapter:in_clk_0_clk, avalon_st_adapter_001:in_clk_0_clk, master_0:clk_clk, mm_interconnect_1:PLL_using_AD1939_MCLK_outclk0_clk, pFIR_Testing_0:clk, rst_controller:clk]
	signal hps_h2f_axi_master_awburst                                    : std_logic_vector(1 downto 0);  -- hps:h2f_AWBURST -> mm_interconnect_0:hps_h2f_axi_master_awburst
	signal hps_h2f_axi_master_arlen                                      : std_logic_vector(3 downto 0);  -- hps:h2f_ARLEN -> mm_interconnect_0:hps_h2f_axi_master_arlen
	signal hps_h2f_axi_master_wstrb                                      : std_logic_vector(7 downto 0);  -- hps:h2f_WSTRB -> mm_interconnect_0:hps_h2f_axi_master_wstrb
	signal hps_h2f_axi_master_wready                                     : std_logic;                     -- mm_interconnect_0:hps_h2f_axi_master_wready -> hps:h2f_WREADY
	signal hps_h2f_axi_master_rid                                        : std_logic_vector(11 downto 0); -- mm_interconnect_0:hps_h2f_axi_master_rid -> hps:h2f_RID
	signal hps_h2f_axi_master_rready                                     : std_logic;                     -- hps:h2f_RREADY -> mm_interconnect_0:hps_h2f_axi_master_rready
	signal hps_h2f_axi_master_awlen                                      : std_logic_vector(3 downto 0);  -- hps:h2f_AWLEN -> mm_interconnect_0:hps_h2f_axi_master_awlen
	signal hps_h2f_axi_master_wid                                        : std_logic_vector(11 downto 0); -- hps:h2f_WID -> mm_interconnect_0:hps_h2f_axi_master_wid
	signal hps_h2f_axi_master_arcache                                    : std_logic_vector(3 downto 0);  -- hps:h2f_ARCACHE -> mm_interconnect_0:hps_h2f_axi_master_arcache
	signal hps_h2f_axi_master_wvalid                                     : std_logic;                     -- hps:h2f_WVALID -> mm_interconnect_0:hps_h2f_axi_master_wvalid
	signal hps_h2f_axi_master_araddr                                     : std_logic_vector(29 downto 0); -- hps:h2f_ARADDR -> mm_interconnect_0:hps_h2f_axi_master_araddr
	signal hps_h2f_axi_master_arprot                                     : std_logic_vector(2 downto 0);  -- hps:h2f_ARPROT -> mm_interconnect_0:hps_h2f_axi_master_arprot
	signal hps_h2f_axi_master_awprot                                     : std_logic_vector(2 downto 0);  -- hps:h2f_AWPROT -> mm_interconnect_0:hps_h2f_axi_master_awprot
	signal hps_h2f_axi_master_wdata                                      : std_logic_vector(63 downto 0); -- hps:h2f_WDATA -> mm_interconnect_0:hps_h2f_axi_master_wdata
	signal hps_h2f_axi_master_arvalid                                    : std_logic;                     -- hps:h2f_ARVALID -> mm_interconnect_0:hps_h2f_axi_master_arvalid
	signal hps_h2f_axi_master_awcache                                    : std_logic_vector(3 downto 0);  -- hps:h2f_AWCACHE -> mm_interconnect_0:hps_h2f_axi_master_awcache
	signal hps_h2f_axi_master_arid                                       : std_logic_vector(11 downto 0); -- hps:h2f_ARID -> mm_interconnect_0:hps_h2f_axi_master_arid
	signal hps_h2f_axi_master_arlock                                     : std_logic_vector(1 downto 0);  -- hps:h2f_ARLOCK -> mm_interconnect_0:hps_h2f_axi_master_arlock
	signal hps_h2f_axi_master_awlock                                     : std_logic_vector(1 downto 0);  -- hps:h2f_AWLOCK -> mm_interconnect_0:hps_h2f_axi_master_awlock
	signal hps_h2f_axi_master_awaddr                                     : std_logic_vector(29 downto 0); -- hps:h2f_AWADDR -> mm_interconnect_0:hps_h2f_axi_master_awaddr
	signal hps_h2f_axi_master_bresp                                      : std_logic_vector(1 downto 0);  -- mm_interconnect_0:hps_h2f_axi_master_bresp -> hps:h2f_BRESP
	signal hps_h2f_axi_master_arready                                    : std_logic;                     -- mm_interconnect_0:hps_h2f_axi_master_arready -> hps:h2f_ARREADY
	signal hps_h2f_axi_master_rdata                                      : std_logic_vector(63 downto 0); -- mm_interconnect_0:hps_h2f_axi_master_rdata -> hps:h2f_RDATA
	signal hps_h2f_axi_master_awready                                    : std_logic;                     -- mm_interconnect_0:hps_h2f_axi_master_awready -> hps:h2f_AWREADY
	signal hps_h2f_axi_master_arburst                                    : std_logic_vector(1 downto 0);  -- hps:h2f_ARBURST -> mm_interconnect_0:hps_h2f_axi_master_arburst
	signal hps_h2f_axi_master_arsize                                     : std_logic_vector(2 downto 0);  -- hps:h2f_ARSIZE -> mm_interconnect_0:hps_h2f_axi_master_arsize
	signal hps_h2f_axi_master_bready                                     : std_logic;                     -- hps:h2f_BREADY -> mm_interconnect_0:hps_h2f_axi_master_bready
	signal hps_h2f_axi_master_rlast                                      : std_logic;                     -- mm_interconnect_0:hps_h2f_axi_master_rlast -> hps:h2f_RLAST
	signal hps_h2f_axi_master_wlast                                      : std_logic;                     -- hps:h2f_WLAST -> mm_interconnect_0:hps_h2f_axi_master_wlast
	signal hps_h2f_axi_master_rresp                                      : std_logic_vector(1 downto 0);  -- mm_interconnect_0:hps_h2f_axi_master_rresp -> hps:h2f_RRESP
	signal hps_h2f_axi_master_awid                                       : std_logic_vector(11 downto 0); -- hps:h2f_AWID -> mm_interconnect_0:hps_h2f_axi_master_awid
	signal hps_h2f_axi_master_bid                                        : std_logic_vector(11 downto 0); -- mm_interconnect_0:hps_h2f_axi_master_bid -> hps:h2f_BID
	signal hps_h2f_axi_master_bvalid                                     : std_logic;                     -- mm_interconnect_0:hps_h2f_axi_master_bvalid -> hps:h2f_BVALID
	signal hps_h2f_axi_master_awsize                                     : std_logic_vector(2 downto 0);  -- hps:h2f_AWSIZE -> mm_interconnect_0:hps_h2f_axi_master_awsize
	signal hps_h2f_axi_master_awvalid                                    : std_logic;                     -- hps:h2f_AWVALID -> mm_interconnect_0:hps_h2f_axi_master_awvalid
	signal hps_h2f_axi_master_rvalid                                     : std_logic;                     -- mm_interconnect_0:hps_h2f_axi_master_rvalid -> hps:h2f_RVALID
	signal mm_interconnect_0_onchip_memory_s1_chipselect                 : std_logic;                     -- mm_interconnect_0:onchip_memory_s1_chipselect -> onchip_memory:chipselect
	signal mm_interconnect_0_onchip_memory_s1_readdata                   : std_logic_vector(63 downto 0); -- onchip_memory:readdata -> mm_interconnect_0:onchip_memory_s1_readdata
	signal mm_interconnect_0_onchip_memory_s1_address                    : std_logic_vector(12 downto 0); -- mm_interconnect_0:onchip_memory_s1_address -> onchip_memory:address
	signal mm_interconnect_0_onchip_memory_s1_byteenable                 : std_logic_vector(7 downto 0);  -- mm_interconnect_0:onchip_memory_s1_byteenable -> onchip_memory:byteenable
	signal mm_interconnect_0_onchip_memory_s1_write                      : std_logic;                     -- mm_interconnect_0:onchip_memory_s1_write -> onchip_memory:write
	signal mm_interconnect_0_onchip_memory_s1_writedata                  : std_logic_vector(63 downto 0); -- mm_interconnect_0:onchip_memory_s1_writedata -> onchip_memory:writedata
	signal mm_interconnect_0_onchip_memory_s1_clken                      : std_logic;                     -- mm_interconnect_0:onchip_memory_s1_clken -> onchip_memory:clken
	signal hps_h2f_lw_axi_master_awburst                                 : std_logic_vector(1 downto 0);  -- hps:h2f_lw_AWBURST -> mm_interconnect_1:hps_h2f_lw_axi_master_awburst
	signal hps_h2f_lw_axi_master_arlen                                   : std_logic_vector(3 downto 0);  -- hps:h2f_lw_ARLEN -> mm_interconnect_1:hps_h2f_lw_axi_master_arlen
	signal hps_h2f_lw_axi_master_wstrb                                   : std_logic_vector(3 downto 0);  -- hps:h2f_lw_WSTRB -> mm_interconnect_1:hps_h2f_lw_axi_master_wstrb
	signal hps_h2f_lw_axi_master_wready                                  : std_logic;                     -- mm_interconnect_1:hps_h2f_lw_axi_master_wready -> hps:h2f_lw_WREADY
	signal hps_h2f_lw_axi_master_rid                                     : std_logic_vector(11 downto 0); -- mm_interconnect_1:hps_h2f_lw_axi_master_rid -> hps:h2f_lw_RID
	signal hps_h2f_lw_axi_master_rready                                  : std_logic;                     -- hps:h2f_lw_RREADY -> mm_interconnect_1:hps_h2f_lw_axi_master_rready
	signal hps_h2f_lw_axi_master_awlen                                   : std_logic_vector(3 downto 0);  -- hps:h2f_lw_AWLEN -> mm_interconnect_1:hps_h2f_lw_axi_master_awlen
	signal hps_h2f_lw_axi_master_wid                                     : std_logic_vector(11 downto 0); -- hps:h2f_lw_WID -> mm_interconnect_1:hps_h2f_lw_axi_master_wid
	signal hps_h2f_lw_axi_master_arcache                                 : std_logic_vector(3 downto 0);  -- hps:h2f_lw_ARCACHE -> mm_interconnect_1:hps_h2f_lw_axi_master_arcache
	signal hps_h2f_lw_axi_master_wvalid                                  : std_logic;                     -- hps:h2f_lw_WVALID -> mm_interconnect_1:hps_h2f_lw_axi_master_wvalid
	signal hps_h2f_lw_axi_master_araddr                                  : std_logic_vector(20 downto 0); -- hps:h2f_lw_ARADDR -> mm_interconnect_1:hps_h2f_lw_axi_master_araddr
	signal hps_h2f_lw_axi_master_arprot                                  : std_logic_vector(2 downto 0);  -- hps:h2f_lw_ARPROT -> mm_interconnect_1:hps_h2f_lw_axi_master_arprot
	signal hps_h2f_lw_axi_master_awprot                                  : std_logic_vector(2 downto 0);  -- hps:h2f_lw_AWPROT -> mm_interconnect_1:hps_h2f_lw_axi_master_awprot
	signal hps_h2f_lw_axi_master_wdata                                   : std_logic_vector(31 downto 0); -- hps:h2f_lw_WDATA -> mm_interconnect_1:hps_h2f_lw_axi_master_wdata
	signal hps_h2f_lw_axi_master_arvalid                                 : std_logic;                     -- hps:h2f_lw_ARVALID -> mm_interconnect_1:hps_h2f_lw_axi_master_arvalid
	signal hps_h2f_lw_axi_master_awcache                                 : std_logic_vector(3 downto 0);  -- hps:h2f_lw_AWCACHE -> mm_interconnect_1:hps_h2f_lw_axi_master_awcache
	signal hps_h2f_lw_axi_master_arid                                    : std_logic_vector(11 downto 0); -- hps:h2f_lw_ARID -> mm_interconnect_1:hps_h2f_lw_axi_master_arid
	signal hps_h2f_lw_axi_master_arlock                                  : std_logic_vector(1 downto 0);  -- hps:h2f_lw_ARLOCK -> mm_interconnect_1:hps_h2f_lw_axi_master_arlock
	signal hps_h2f_lw_axi_master_awlock                                  : std_logic_vector(1 downto 0);  -- hps:h2f_lw_AWLOCK -> mm_interconnect_1:hps_h2f_lw_axi_master_awlock
	signal hps_h2f_lw_axi_master_awaddr                                  : std_logic_vector(20 downto 0); -- hps:h2f_lw_AWADDR -> mm_interconnect_1:hps_h2f_lw_axi_master_awaddr
	signal hps_h2f_lw_axi_master_bresp                                   : std_logic_vector(1 downto 0);  -- mm_interconnect_1:hps_h2f_lw_axi_master_bresp -> hps:h2f_lw_BRESP
	signal hps_h2f_lw_axi_master_arready                                 : std_logic;                     -- mm_interconnect_1:hps_h2f_lw_axi_master_arready -> hps:h2f_lw_ARREADY
	signal hps_h2f_lw_axi_master_rdata                                   : std_logic_vector(31 downto 0); -- mm_interconnect_1:hps_h2f_lw_axi_master_rdata -> hps:h2f_lw_RDATA
	signal hps_h2f_lw_axi_master_awready                                 : std_logic;                     -- mm_interconnect_1:hps_h2f_lw_axi_master_awready -> hps:h2f_lw_AWREADY
	signal hps_h2f_lw_axi_master_arburst                                 : std_logic_vector(1 downto 0);  -- hps:h2f_lw_ARBURST -> mm_interconnect_1:hps_h2f_lw_axi_master_arburst
	signal hps_h2f_lw_axi_master_arsize                                  : std_logic_vector(2 downto 0);  -- hps:h2f_lw_ARSIZE -> mm_interconnect_1:hps_h2f_lw_axi_master_arsize
	signal hps_h2f_lw_axi_master_bready                                  : std_logic;                     -- hps:h2f_lw_BREADY -> mm_interconnect_1:hps_h2f_lw_axi_master_bready
	signal hps_h2f_lw_axi_master_rlast                                   : std_logic;                     -- mm_interconnect_1:hps_h2f_lw_axi_master_rlast -> hps:h2f_lw_RLAST
	signal hps_h2f_lw_axi_master_wlast                                   : std_logic;                     -- hps:h2f_lw_WLAST -> mm_interconnect_1:hps_h2f_lw_axi_master_wlast
	signal hps_h2f_lw_axi_master_rresp                                   : std_logic_vector(1 downto 0);  -- mm_interconnect_1:hps_h2f_lw_axi_master_rresp -> hps:h2f_lw_RRESP
	signal hps_h2f_lw_axi_master_awid                                    : std_logic_vector(11 downto 0); -- hps:h2f_lw_AWID -> mm_interconnect_1:hps_h2f_lw_axi_master_awid
	signal hps_h2f_lw_axi_master_bid                                     : std_logic_vector(11 downto 0); -- mm_interconnect_1:hps_h2f_lw_axi_master_bid -> hps:h2f_lw_BID
	signal hps_h2f_lw_axi_master_bvalid                                  : std_logic;                     -- mm_interconnect_1:hps_h2f_lw_axi_master_bvalid -> hps:h2f_lw_BVALID
	signal hps_h2f_lw_axi_master_awsize                                  : std_logic_vector(2 downto 0);  -- hps:h2f_lw_AWSIZE -> mm_interconnect_1:hps_h2f_lw_axi_master_awsize
	signal hps_h2f_lw_axi_master_awvalid                                 : std_logic;                     -- hps:h2f_lw_AWVALID -> mm_interconnect_1:hps_h2f_lw_axi_master_awvalid
	signal hps_h2f_lw_axi_master_rvalid                                  : std_logic;                     -- mm_interconnect_1:hps_h2f_lw_axi_master_rvalid -> hps:h2f_lw_RVALID
	signal master_0_master_readdata                                      : std_logic_vector(31 downto 0); -- mm_interconnect_1:master_0_master_readdata -> master_0:master_readdata
	signal master_0_master_waitrequest                                   : std_logic;                     -- mm_interconnect_1:master_0_master_waitrequest -> master_0:master_waitrequest
	signal master_0_master_address                                       : std_logic_vector(31 downto 0); -- master_0:master_address -> mm_interconnect_1:master_0_master_address
	signal master_0_master_read                                          : std_logic;                     -- master_0:master_read -> mm_interconnect_1:master_0_master_read
	signal master_0_master_byteenable                                    : std_logic_vector(3 downto 0);  -- master_0:master_byteenable -> mm_interconnect_1:master_0_master_byteenable
	signal master_0_master_readdatavalid                                 : std_logic;                     -- mm_interconnect_1:master_0_master_readdatavalid -> master_0:master_readdatavalid
	signal master_0_master_write                                         : std_logic;                     -- master_0:master_write -> mm_interconnect_1:master_0_master_write
	signal master_0_master_writedata                                     : std_logic_vector(31 downto 0); -- master_0:master_writedata -> mm_interconnect_1:master_0_master_writedata
	signal mm_interconnect_1_jtag_uart_avalon_jtag_slave_chipselect      : std_logic;                     -- mm_interconnect_1:jtag_uart_avalon_jtag_slave_chipselect -> jtag_uart:av_chipselect
	signal mm_interconnect_1_jtag_uart_avalon_jtag_slave_readdata        : std_logic_vector(31 downto 0); -- jtag_uart:av_readdata -> mm_interconnect_1:jtag_uart_avalon_jtag_slave_readdata
	signal mm_interconnect_1_jtag_uart_avalon_jtag_slave_waitrequest     : std_logic;                     -- jtag_uart:av_waitrequest -> mm_interconnect_1:jtag_uart_avalon_jtag_slave_waitrequest
	signal mm_interconnect_1_jtag_uart_avalon_jtag_slave_address         : std_logic_vector(0 downto 0);  -- mm_interconnect_1:jtag_uart_avalon_jtag_slave_address -> jtag_uart:av_address
	signal mm_interconnect_1_jtag_uart_avalon_jtag_slave_read            : std_logic;                     -- mm_interconnect_1:jtag_uart_avalon_jtag_slave_read -> mm_interconnect_1_jtag_uart_avalon_jtag_slave_read:in
	signal mm_interconnect_1_jtag_uart_avalon_jtag_slave_write           : std_logic;                     -- mm_interconnect_1:jtag_uart_avalon_jtag_slave_write -> mm_interconnect_1_jtag_uart_avalon_jtag_slave_write:in
	signal mm_interconnect_1_jtag_uart_avalon_jtag_slave_writedata       : std_logic_vector(31 downto 0); -- mm_interconnect_1:jtag_uart_avalon_jtag_slave_writedata -> jtag_uart:av_writedata
	signal mm_interconnect_1_pfir_testing_0_avalon_slave_0_readdata      : std_logic_vector(31 downto 0); -- pFIR_Testing_0:avalon_slave_0_readdata -> mm_interconnect_1:pFIR_Testing_0_avalon_slave_0_readdata
	signal mm_interconnect_1_pfir_testing_0_avalon_slave_0_address       : std_logic_vector(0 downto 0);  -- mm_interconnect_1:pFIR_Testing_0_avalon_slave_0_address -> pFIR_Testing_0:avalon_slave_0_address
	signal mm_interconnect_1_pfir_testing_0_avalon_slave_0_read          : std_logic;                     -- mm_interconnect_1:pFIR_Testing_0_avalon_slave_0_read -> pFIR_Testing_0:avalon_slave_0_read
	signal mm_interconnect_1_pfir_testing_0_avalon_slave_0_write         : std_logic;                     -- mm_interconnect_1:pFIR_Testing_0_avalon_slave_0_write -> pFIR_Testing_0:avalon_slave_0_write
	signal mm_interconnect_1_pfir_testing_0_avalon_slave_0_writedata     : std_logic_vector(31 downto 0); -- mm_interconnect_1:pFIR_Testing_0_avalon_slave_0_writedata -> pFIR_Testing_0:avalon_slave_0_writedata
	signal mm_interconnect_1_pfir_testing_0_avalon_slave_1_readdata      : std_logic_vector(31 downto 0); -- pFIR_Testing_0:avalon_slave_1_readdata -> mm_interconnect_1:pFIR_Testing_0_avalon_slave_1_readdata
	signal mm_interconnect_1_pfir_testing_0_avalon_slave_1_address       : std_logic_vector(8 downto 0);  -- mm_interconnect_1:pFIR_Testing_0_avalon_slave_1_address -> pFIR_Testing_0:avalon_slave_1_address
	signal mm_interconnect_1_pfir_testing_0_avalon_slave_1_read          : std_logic;                     -- mm_interconnect_1:pFIR_Testing_0_avalon_slave_1_read -> pFIR_Testing_0:avalon_slave_1_read
	signal mm_interconnect_1_pfir_testing_0_avalon_slave_1_write         : std_logic;                     -- mm_interconnect_1:pFIR_Testing_0_avalon_slave_1_write -> pFIR_Testing_0:avalon_slave_1_write
	signal mm_interconnect_1_pfir_testing_0_avalon_slave_1_writedata     : std_logic_vector(31 downto 0); -- mm_interconnect_1:pFIR_Testing_0_avalon_slave_1_writedata -> pFIR_Testing_0:avalon_slave_1_writedata
	signal mm_interconnect_1_systemid_control_slave_readdata             : std_logic_vector(31 downto 0); -- SystemID:readdata -> mm_interconnect_1:SystemID_control_slave_readdata
	signal mm_interconnect_1_systemid_control_slave_address              : std_logic_vector(0 downto 0);  -- mm_interconnect_1:SystemID_control_slave_address -> SystemID:address
	signal irq_mapper_receiver0_irq                                      : std_logic;                     -- jtag_uart:av_irq -> irq_mapper:receiver0_irq
	signal hps_f2h_irq0_irq                                              : std_logic_vector(31 downto 0); -- irq_mapper:sender_irq -> hps:f2h_irq_p0
	signal hps_f2h_irq1_irq                                              : std_logic_vector(31 downto 0); -- irq_mapper_001:sender_irq -> hps:f2h_irq_p1
	signal fe_qsys_ad1939_audio_mini_v1_0_line_in_valid                  : std_logic;                     -- FE_Qsys_AD1939_Audio_Mini_v1_0:AD1939_ADC_valid -> avalon_st_adapter:in_0_valid
	signal fe_qsys_ad1939_audio_mini_v1_0_line_in_data                   : std_logic_vector(31 downto 0); -- FE_Qsys_AD1939_Audio_Mini_v1_0:AD1939_ADC_data -> avalon_st_adapter:in_0_data
	signal fe_qsys_ad1939_audio_mini_v1_0_line_in_channel                : std_logic_vector(1 downto 0);  -- FE_Qsys_AD1939_Audio_Mini_v1_0:AD1939_ADC_channel -> avalon_st_adapter:in_0_channel
	signal fe_qsys_ad1939_audio_mini_v1_0_line_in_error                  : std_logic_vector(1 downto 0);  -- FE_Qsys_AD1939_Audio_Mini_v1_0:AD1939_ADC_error -> avalon_st_adapter:in_0_error
	signal avalon_st_adapter_out_0_valid                                 : std_logic;                     -- avalon_st_adapter:out_0_valid -> pFIR_Testing_0:avalon_sink_valid
	signal avalon_st_adapter_out_0_data                                  : std_logic_vector(31 downto 0); -- avalon_st_adapter:out_0_data -> pFIR_Testing_0:avalon_sink_data
	signal avalon_st_adapter_out_0_channel                               : std_logic_vector(1 downto 0);  -- avalon_st_adapter:out_0_channel -> pFIR_Testing_0:avalon_sink_channel
	signal avalon_st_adapter_out_0_error                                 : std_logic_vector(1 downto 0);  -- avalon_st_adapter:out_0_error -> pFIR_Testing_0:avalon_sink_error
	signal pfir_testing_0_avalon_streaming_source_valid                  : std_logic;                     -- pFIR_Testing_0:avalon_source_valid -> avalon_st_adapter_001:in_0_valid
	signal pfir_testing_0_avalon_streaming_source_data                   : std_logic_vector(31 downto 0); -- pFIR_Testing_0:avalon_source_data -> avalon_st_adapter_001:in_0_data
	signal pfir_testing_0_avalon_streaming_source_channel                : std_logic_vector(1 downto 0);  -- pFIR_Testing_0:avalon_source_channel -> avalon_st_adapter_001:in_0_channel
	signal pfir_testing_0_avalon_streaming_source_error                  : std_logic_vector(1 downto 0);  -- pFIR_Testing_0:avalon_source_error -> avalon_st_adapter_001:in_0_error
	signal avalon_st_adapter_001_out_0_valid                             : std_logic;                     -- avalon_st_adapter_001:out_0_valid -> FE_Qsys_AD1939_Audio_Mini_v1_0:AD1939_DAC_valid
	signal avalon_st_adapter_001_out_0_data                              : std_logic_vector(31 downto 0); -- avalon_st_adapter_001:out_0_data -> FE_Qsys_AD1939_Audio_Mini_v1_0:AD1939_DAC_data
	signal avalon_st_adapter_001_out_0_channel                           : std_logic_vector(1 downto 0);  -- avalon_st_adapter_001:out_0_channel -> FE_Qsys_AD1939_Audio_Mini_v1_0:AD1939_DAC_channel
	signal avalon_st_adapter_001_out_0_error                             : std_logic_vector(1 downto 0);  -- avalon_st_adapter_001:out_0_error -> FE_Qsys_AD1939_Audio_Mini_v1_0:AD1939_DAC_error
	signal rst_controller_reset_out_reset                                : std_logic;                     -- rst_controller:reset_out -> [FE_Qsys_AD1939_Audio_Mini_v1_0:sys_reset, avalon_st_adapter:in_rst_0_reset, avalon_st_adapter_001:in_rst_0_reset, mm_interconnect_1:master_0_clk_reset_reset_bridge_in_reset_reset, mm_interconnect_1:pFIR_Testing_0_reset_reset_bridge_in_reset_reset, pFIR_Testing_0:reset]
	signal rst_controller_001_reset_out_reset                            : std_logic;                     -- rst_controller_001:reset_out -> [mm_interconnect_0:onchip_memory_reset1_reset_bridge_in_reset_reset, mm_interconnect_1:SystemID_reset_reset_bridge_in_reset_reset, onchip_memory:reset, rst_controller_001_reset_out_reset:in, rst_translator:in_reset]
	signal rst_controller_001_reset_out_reset_req                        : std_logic;                     -- rst_controller_001:reset_req -> [onchip_memory:reset_req, rst_translator:reset_req_in]
	signal rst_controller_002_reset_out_reset                            : std_logic;                     -- rst_controller_002:reset_out -> [mm_interconnect_1:jtag_uart_reset_reset_bridge_in_reset_reset, rst_controller_002_reset_out_reset:in]
	signal master_0_master_reset_reset                                   : std_logic;                     -- master_0:master_reset_reset -> rst_controller_002:reset_in1
	signal rst_controller_003_reset_out_reset                            : std_logic;                     -- rst_controller_003:reset_out -> [mm_interconnect_0:hps_h2f_axi_master_agent_clk_reset_reset_bridge_in_reset_reset, mm_interconnect_1:hps_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset_reset]
	signal hps_h2f_reset_reset_n_ports_inv                               : std_logic;                     -- hps_h2f_reset_reset_n:inv -> rst_controller_003:reset_in0
	signal reset_reset_n_ports_inv                                       : std_logic;                     -- reset_reset_n:inv -> [PLL_using_AD1939_MCLK:rst, master_0:clk_reset_reset, rst_controller:reset_in0, rst_controller_001:reset_in0, rst_controller_002:reset_in0]
	signal mm_interconnect_1_jtag_uart_avalon_jtag_slave_read_ports_inv  : std_logic;                     -- mm_interconnect_1_jtag_uart_avalon_jtag_slave_read:inv -> jtag_uart:av_read_n
	signal mm_interconnect_1_jtag_uart_avalon_jtag_slave_write_ports_inv : std_logic;                     -- mm_interconnect_1_jtag_uart_avalon_jtag_slave_write:inv -> jtag_uart:av_write_n
	signal rst_controller_001_reset_out_reset_ports_inv                  : std_logic;                     -- rst_controller_001_reset_out_reset:inv -> SystemID:reset_n
	signal rst_controller_002_reset_out_reset_ports_inv                  : std_logic;                     -- rst_controller_002_reset_out_reset:inv -> jtag_uart:rst_n

begin

	fe_qsys_ad1939_audio_mini_v1_0 : component AD1939_hps_audio_mini
		port map (
			sys_clk            => pll_using_ad1939_mclk_outclk0_clk,              --           sys_clk.clk
			sys_reset          => rst_controller_reset_out_reset,                 --         sys_reset.reset
			AD1939_ADC_ABCLK   => ad1939_abclk_clk,                               --         clk_abclk.clk
			AD1939_ADC_ALRCLK  => ad1939_alrclk_clk,                              --        clk_alrclk.clk
			AD1939_ADC_channel => fe_qsys_ad1939_audio_mini_v1_0_line_in_channel, --           Line_In.channel
			AD1939_ADC_data    => fe_qsys_ad1939_audio_mini_v1_0_line_in_data,    --                  .data
			AD1939_ADC_error   => fe_qsys_ad1939_audio_mini_v1_0_line_in_error,   --                  .error
			AD1939_ADC_valid   => fe_qsys_ad1939_audio_mini_v1_0_line_in_valid,   --                  .valid
			AD1939_DAC_channel => avalon_st_adapter_001_out_0_channel,            --     Headphone_Out.channel
			AD1939_DAC_data    => avalon_st_adapter_001_out_0_data,               --                  .data
			AD1939_DAC_error   => avalon_st_adapter_001_out_0_error,              --                  .error
			AD1939_DAC_valid   => avalon_st_adapter_001_out_0_valid,              --                  .valid
			AD1939_ADC_ASDATA2 => ad1939_physical_asdata2,                        -- connect_to_AD1939.asdata2
			AD1939_DAC_DBCLK   => ad1939_physical_dbclk,                          --                  .dbclk
			AD1939_DAC_DLRCLK  => ad1939_physical_dlrclk,                         --                  .dlrclk
			AD1939_DAC_DSDATA1 => ad1939_physical_dsdata1                         --                  .dsdata1
		);

	pll_using_ad1939_mclk : component soc_system_PLL_using_AD1939_MCLK
		port map (
			refclk   => ad1939_mclk_clk,                   --  refclk.clk
			rst      => reset_reset_n_ports_inv,           --   reset.reset
			outclk_0 => pll_using_ad1939_mclk_outclk0_clk, -- outclk0.clk
			locked   => open                               -- (terminated)
		);

	systemid : component soc_system_SystemID
		port map (
			clock    => clk_clk,                                             --           clk.clk
			reset_n  => rst_controller_001_reset_out_reset_ports_inv,        --         reset.reset_n
			readdata => mm_interconnect_1_systemid_control_slave_readdata,   -- control_slave.readdata
			address  => mm_interconnect_1_systemid_control_slave_address(0)  --              .address
		);

	hps : component soc_system_hps
		generic map (
			F2S_Width => 3,
			S2F_Width => 2
		)
		port map (
			h2f_cold_rst_n           => open,                                --      h2f_cold_reset.reset_n
			f2h_cold_rst_req_n       => hps_f2h_cold_reset_req_reset_n,      --  f2h_cold_reset_req.reset_n
			f2h_dbg_rst_req_n        => hps_f2h_debug_reset_req_reset_n,     -- f2h_debug_reset_req.reset_n
			f2h_warm_rst_req_n       => hps_f2h_warm_reset_req_reset_n,      --  f2h_warm_reset_req.reset_n
			spim0_txd                => hps_spim0_txd,                       --               spim0.txd
			spim0_rxd                => hps_spim0_rxd,                       --                    .rxd
			spim0_ss_in_n            => hps_spim0_ss_in_n,                   --                    .ss_in_n
			spim0_ssi_oe_n           => hps_spim0_ssi_oe_n,                  --                    .ssi_oe_n
			spim0_ss_0_n             => hps_spim0_ss_0_n,                    --                    .ss_0_n
			spim0_ss_1_n             => hps_spim0_ss_1_n,                    --                    .ss_1_n
			spim0_ss_2_n             => hps_spim0_ss_2_n,                    --                    .ss_2_n
			spim0_ss_3_n             => hps_spim0_ss_3_n,                    --                    .ss_3_n
			spim0_sclk_out           => hps_spim0_sclk_out_clk,              --      spim0_sclk_out.clk
			i2c0_scl                 => hps_i2c0_scl_in_clk,                 --         i2c0_scl_in.clk
			i2c0_out_clk             => hps_i2c0_clk_clk,                    --            i2c0_clk.clk
			i2c0_out_data            => hps_i2c0_out_data,                   --                i2c0.out_data
			i2c0_sda                 => hps_i2c0_sda,                        --                    .sda
			mem_a                    => memory_mem_a,                        --              memory.mem_a
			mem_ba                   => memory_mem_ba,                       --                    .mem_ba
			mem_ck                   => memory_mem_ck,                       --                    .mem_ck
			mem_ck_n                 => memory_mem_ck_n,                     --                    .mem_ck_n
			mem_cke                  => memory_mem_cke,                      --                    .mem_cke
			mem_cs_n                 => memory_mem_cs_n,                     --                    .mem_cs_n
			mem_ras_n                => memory_mem_ras_n,                    --                    .mem_ras_n
			mem_cas_n                => memory_mem_cas_n,                    --                    .mem_cas_n
			mem_we_n                 => memory_mem_we_n,                     --                    .mem_we_n
			mem_reset_n              => memory_mem_reset_n,                  --                    .mem_reset_n
			mem_dq                   => memory_mem_dq,                       --                    .mem_dq
			mem_dqs                  => memory_mem_dqs,                      --                    .mem_dqs
			mem_dqs_n                => memory_mem_dqs_n,                    --                    .mem_dqs_n
			mem_odt                  => memory_mem_odt,                      --                    .mem_odt
			mem_dm                   => memory_mem_dm,                       --                    .mem_dm
			oct_rzqin                => memory_oct_rzqin,                    --                    .oct_rzqin
			hps_io_emac1_inst_TX_CLK => hps_hps_io_hps_io_emac1_inst_TX_CLK, --              hps_io.hps_io_emac1_inst_TX_CLK
			hps_io_emac1_inst_TXD0   => hps_hps_io_hps_io_emac1_inst_TXD0,   --                    .hps_io_emac1_inst_TXD0
			hps_io_emac1_inst_TXD1   => hps_hps_io_hps_io_emac1_inst_TXD1,   --                    .hps_io_emac1_inst_TXD1
			hps_io_emac1_inst_TXD2   => hps_hps_io_hps_io_emac1_inst_TXD2,   --                    .hps_io_emac1_inst_TXD2
			hps_io_emac1_inst_TXD3   => hps_hps_io_hps_io_emac1_inst_TXD3,   --                    .hps_io_emac1_inst_TXD3
			hps_io_emac1_inst_RXD0   => hps_hps_io_hps_io_emac1_inst_RXD0,   --                    .hps_io_emac1_inst_RXD0
			hps_io_emac1_inst_MDIO   => hps_hps_io_hps_io_emac1_inst_MDIO,   --                    .hps_io_emac1_inst_MDIO
			hps_io_emac1_inst_MDC    => hps_hps_io_hps_io_emac1_inst_MDC,    --                    .hps_io_emac1_inst_MDC
			hps_io_emac1_inst_RX_CTL => hps_hps_io_hps_io_emac1_inst_RX_CTL, --                    .hps_io_emac1_inst_RX_CTL
			hps_io_emac1_inst_TX_CTL => hps_hps_io_hps_io_emac1_inst_TX_CTL, --                    .hps_io_emac1_inst_TX_CTL
			hps_io_emac1_inst_RX_CLK => hps_hps_io_hps_io_emac1_inst_RX_CLK, --                    .hps_io_emac1_inst_RX_CLK
			hps_io_emac1_inst_RXD1   => hps_hps_io_hps_io_emac1_inst_RXD1,   --                    .hps_io_emac1_inst_RXD1
			hps_io_emac1_inst_RXD2   => hps_hps_io_hps_io_emac1_inst_RXD2,   --                    .hps_io_emac1_inst_RXD2
			hps_io_emac1_inst_RXD3   => hps_hps_io_hps_io_emac1_inst_RXD3,   --                    .hps_io_emac1_inst_RXD3
			hps_io_sdio_inst_CMD     => hps_hps_io_hps_io_sdio_inst_CMD,     --                    .hps_io_sdio_inst_CMD
			hps_io_sdio_inst_D0      => hps_hps_io_hps_io_sdio_inst_D0,      --                    .hps_io_sdio_inst_D0
			hps_io_sdio_inst_D1      => hps_hps_io_hps_io_sdio_inst_D1,      --                    .hps_io_sdio_inst_D1
			hps_io_sdio_inst_CLK     => hps_hps_io_hps_io_sdio_inst_CLK,     --                    .hps_io_sdio_inst_CLK
			hps_io_sdio_inst_D2      => hps_hps_io_hps_io_sdio_inst_D2,      --                    .hps_io_sdio_inst_D2
			hps_io_sdio_inst_D3      => hps_hps_io_hps_io_sdio_inst_D3,      --                    .hps_io_sdio_inst_D3
			hps_io_usb1_inst_D0      => hps_hps_io_hps_io_usb1_inst_D0,      --                    .hps_io_usb1_inst_D0
			hps_io_usb1_inst_D1      => hps_hps_io_hps_io_usb1_inst_D1,      --                    .hps_io_usb1_inst_D1
			hps_io_usb1_inst_D2      => hps_hps_io_hps_io_usb1_inst_D2,      --                    .hps_io_usb1_inst_D2
			hps_io_usb1_inst_D3      => hps_hps_io_hps_io_usb1_inst_D3,      --                    .hps_io_usb1_inst_D3
			hps_io_usb1_inst_D4      => hps_hps_io_hps_io_usb1_inst_D4,      --                    .hps_io_usb1_inst_D4
			hps_io_usb1_inst_D5      => hps_hps_io_hps_io_usb1_inst_D5,      --                    .hps_io_usb1_inst_D5
			hps_io_usb1_inst_D6      => hps_hps_io_hps_io_usb1_inst_D6,      --                    .hps_io_usb1_inst_D6
			hps_io_usb1_inst_D7      => hps_hps_io_hps_io_usb1_inst_D7,      --                    .hps_io_usb1_inst_D7
			hps_io_usb1_inst_CLK     => hps_hps_io_hps_io_usb1_inst_CLK,     --                    .hps_io_usb1_inst_CLK
			hps_io_usb1_inst_STP     => hps_hps_io_hps_io_usb1_inst_STP,     --                    .hps_io_usb1_inst_STP
			hps_io_usb1_inst_DIR     => hps_hps_io_hps_io_usb1_inst_DIR,     --                    .hps_io_usb1_inst_DIR
			hps_io_usb1_inst_NXT     => hps_hps_io_hps_io_usb1_inst_NXT,     --                    .hps_io_usb1_inst_NXT
			hps_io_spim1_inst_CLK    => hps_hps_io_hps_io_spim1_inst_CLK,    --                    .hps_io_spim1_inst_CLK
			hps_io_spim1_inst_MOSI   => hps_hps_io_hps_io_spim1_inst_MOSI,   --                    .hps_io_spim1_inst_MOSI
			hps_io_spim1_inst_MISO   => hps_hps_io_hps_io_spim1_inst_MISO,   --                    .hps_io_spim1_inst_MISO
			hps_io_spim1_inst_SS0    => hps_hps_io_hps_io_spim1_inst_SS0,    --                    .hps_io_spim1_inst_SS0
			hps_io_uart0_inst_RX     => hps_hps_io_hps_io_uart0_inst_RX,     --                    .hps_io_uart0_inst_RX
			hps_io_uart0_inst_TX     => hps_hps_io_hps_io_uart0_inst_TX,     --                    .hps_io_uart0_inst_TX
			hps_io_i2c1_inst_SDA     => hps_hps_io_hps_io_i2c1_inst_SDA,     --                    .hps_io_i2c1_inst_SDA
			hps_io_i2c1_inst_SCL     => hps_hps_io_hps_io_i2c1_inst_SCL,     --                    .hps_io_i2c1_inst_SCL
			hps_io_gpio_inst_GPIO09  => hps_hps_io_hps_io_gpio_inst_GPIO09,  --                    .hps_io_gpio_inst_GPIO09
			hps_io_gpio_inst_GPIO35  => hps_hps_io_hps_io_gpio_inst_GPIO35,  --                    .hps_io_gpio_inst_GPIO35
			hps_io_gpio_inst_GPIO40  => hps_hps_io_hps_io_gpio_inst_GPIO40,  --                    .hps_io_gpio_inst_GPIO40
			hps_io_gpio_inst_GPIO53  => hps_hps_io_hps_io_gpio_inst_GPIO53,  --                    .hps_io_gpio_inst_GPIO53
			hps_io_gpio_inst_GPIO54  => hps_hps_io_hps_io_gpio_inst_GPIO54,  --                    .hps_io_gpio_inst_GPIO54
			hps_io_gpio_inst_GPIO61  => hps_hps_io_hps_io_gpio_inst_GPIO61,  --                    .hps_io_gpio_inst_GPIO61
			h2f_rst_n                => hps_h2f_reset_reset,                 --           h2f_reset.reset_n
			h2f_axi_clk              => clk_clk,                             --       h2f_axi_clock.clk
			h2f_AWID                 => hps_h2f_axi_master_awid,             --      h2f_axi_master.awid
			h2f_AWADDR               => hps_h2f_axi_master_awaddr,           --                    .awaddr
			h2f_AWLEN                => hps_h2f_axi_master_awlen,            --                    .awlen
			h2f_AWSIZE               => hps_h2f_axi_master_awsize,           --                    .awsize
			h2f_AWBURST              => hps_h2f_axi_master_awburst,          --                    .awburst
			h2f_AWLOCK               => hps_h2f_axi_master_awlock,           --                    .awlock
			h2f_AWCACHE              => hps_h2f_axi_master_awcache,          --                    .awcache
			h2f_AWPROT               => hps_h2f_axi_master_awprot,           --                    .awprot
			h2f_AWVALID              => hps_h2f_axi_master_awvalid,          --                    .awvalid
			h2f_AWREADY              => hps_h2f_axi_master_awready,          --                    .awready
			h2f_WID                  => hps_h2f_axi_master_wid,              --                    .wid
			h2f_WDATA                => hps_h2f_axi_master_wdata,            --                    .wdata
			h2f_WSTRB                => hps_h2f_axi_master_wstrb,            --                    .wstrb
			h2f_WLAST                => hps_h2f_axi_master_wlast,            --                    .wlast
			h2f_WVALID               => hps_h2f_axi_master_wvalid,           --                    .wvalid
			h2f_WREADY               => hps_h2f_axi_master_wready,           --                    .wready
			h2f_BID                  => hps_h2f_axi_master_bid,              --                    .bid
			h2f_BRESP                => hps_h2f_axi_master_bresp,            --                    .bresp
			h2f_BVALID               => hps_h2f_axi_master_bvalid,           --                    .bvalid
			h2f_BREADY               => hps_h2f_axi_master_bready,           --                    .bready
			h2f_ARID                 => hps_h2f_axi_master_arid,             --                    .arid
			h2f_ARADDR               => hps_h2f_axi_master_araddr,           --                    .araddr
			h2f_ARLEN                => hps_h2f_axi_master_arlen,            --                    .arlen
			h2f_ARSIZE               => hps_h2f_axi_master_arsize,           --                    .arsize
			h2f_ARBURST              => hps_h2f_axi_master_arburst,          --                    .arburst
			h2f_ARLOCK               => hps_h2f_axi_master_arlock,           --                    .arlock
			h2f_ARCACHE              => hps_h2f_axi_master_arcache,          --                    .arcache
			h2f_ARPROT               => hps_h2f_axi_master_arprot,           --                    .arprot
			h2f_ARVALID              => hps_h2f_axi_master_arvalid,          --                    .arvalid
			h2f_ARREADY              => hps_h2f_axi_master_arready,          --                    .arready
			h2f_RID                  => hps_h2f_axi_master_rid,              --                    .rid
			h2f_RDATA                => hps_h2f_axi_master_rdata,            --                    .rdata
			h2f_RRESP                => hps_h2f_axi_master_rresp,            --                    .rresp
			h2f_RLAST                => hps_h2f_axi_master_rlast,            --                    .rlast
			h2f_RVALID               => hps_h2f_axi_master_rvalid,           --                    .rvalid
			h2f_RREADY               => hps_h2f_axi_master_rready,           --                    .rready
			f2h_axi_clk              => clk_clk,                             --       f2h_axi_clock.clk
			f2h_AWID                 => open,                                --       f2h_axi_slave.awid
			f2h_AWADDR               => open,                                --                    .awaddr
			f2h_AWLEN                => open,                                --                    .awlen
			f2h_AWSIZE               => open,                                --                    .awsize
			f2h_AWBURST              => open,                                --                    .awburst
			f2h_AWLOCK               => open,                                --                    .awlock
			f2h_AWCACHE              => open,                                --                    .awcache
			f2h_AWPROT               => open,                                --                    .awprot
			f2h_AWVALID              => open,                                --                    .awvalid
			f2h_AWREADY              => open,                                --                    .awready
			f2h_AWUSER               => open,                                --                    .awuser
			f2h_WID                  => open,                                --                    .wid
			f2h_WDATA                => open,                                --                    .wdata
			f2h_WSTRB                => open,                                --                    .wstrb
			f2h_WLAST                => open,                                --                    .wlast
			f2h_WVALID               => open,                                --                    .wvalid
			f2h_WREADY               => open,                                --                    .wready
			f2h_BID                  => open,                                --                    .bid
			f2h_BRESP                => open,                                --                    .bresp
			f2h_BVALID               => open,                                --                    .bvalid
			f2h_BREADY               => open,                                --                    .bready
			f2h_ARID                 => open,                                --                    .arid
			f2h_ARADDR               => open,                                --                    .araddr
			f2h_ARLEN                => open,                                --                    .arlen
			f2h_ARSIZE               => open,                                --                    .arsize
			f2h_ARBURST              => open,                                --                    .arburst
			f2h_ARLOCK               => open,                                --                    .arlock
			f2h_ARCACHE              => open,                                --                    .arcache
			f2h_ARPROT               => open,                                --                    .arprot
			f2h_ARVALID              => open,                                --                    .arvalid
			f2h_ARREADY              => open,                                --                    .arready
			f2h_ARUSER               => open,                                --                    .aruser
			f2h_RID                  => open,                                --                    .rid
			f2h_RDATA                => open,                                --                    .rdata
			f2h_RRESP                => open,                                --                    .rresp
			f2h_RLAST                => open,                                --                    .rlast
			f2h_RVALID               => open,                                --                    .rvalid
			f2h_RREADY               => open,                                --                    .rready
			h2f_lw_axi_clk           => clk_clk,                             --    h2f_lw_axi_clock.clk
			h2f_lw_AWID              => hps_h2f_lw_axi_master_awid,          --   h2f_lw_axi_master.awid
			h2f_lw_AWADDR            => hps_h2f_lw_axi_master_awaddr,        --                    .awaddr
			h2f_lw_AWLEN             => hps_h2f_lw_axi_master_awlen,         --                    .awlen
			h2f_lw_AWSIZE            => hps_h2f_lw_axi_master_awsize,        --                    .awsize
			h2f_lw_AWBURST           => hps_h2f_lw_axi_master_awburst,       --                    .awburst
			h2f_lw_AWLOCK            => hps_h2f_lw_axi_master_awlock,        --                    .awlock
			h2f_lw_AWCACHE           => hps_h2f_lw_axi_master_awcache,       --                    .awcache
			h2f_lw_AWPROT            => hps_h2f_lw_axi_master_awprot,        --                    .awprot
			h2f_lw_AWVALID           => hps_h2f_lw_axi_master_awvalid,       --                    .awvalid
			h2f_lw_AWREADY           => hps_h2f_lw_axi_master_awready,       --                    .awready
			h2f_lw_WID               => hps_h2f_lw_axi_master_wid,           --                    .wid
			h2f_lw_WDATA             => hps_h2f_lw_axi_master_wdata,         --                    .wdata
			h2f_lw_WSTRB             => hps_h2f_lw_axi_master_wstrb,         --                    .wstrb
			h2f_lw_WLAST             => hps_h2f_lw_axi_master_wlast,         --                    .wlast
			h2f_lw_WVALID            => hps_h2f_lw_axi_master_wvalid,        --                    .wvalid
			h2f_lw_WREADY            => hps_h2f_lw_axi_master_wready,        --                    .wready
			h2f_lw_BID               => hps_h2f_lw_axi_master_bid,           --                    .bid
			h2f_lw_BRESP             => hps_h2f_lw_axi_master_bresp,         --                    .bresp
			h2f_lw_BVALID            => hps_h2f_lw_axi_master_bvalid,        --                    .bvalid
			h2f_lw_BREADY            => hps_h2f_lw_axi_master_bready,        --                    .bready
			h2f_lw_ARID              => hps_h2f_lw_axi_master_arid,          --                    .arid
			h2f_lw_ARADDR            => hps_h2f_lw_axi_master_araddr,        --                    .araddr
			h2f_lw_ARLEN             => hps_h2f_lw_axi_master_arlen,         --                    .arlen
			h2f_lw_ARSIZE            => hps_h2f_lw_axi_master_arsize,        --                    .arsize
			h2f_lw_ARBURST           => hps_h2f_lw_axi_master_arburst,       --                    .arburst
			h2f_lw_ARLOCK            => hps_h2f_lw_axi_master_arlock,        --                    .arlock
			h2f_lw_ARCACHE           => hps_h2f_lw_axi_master_arcache,       --                    .arcache
			h2f_lw_ARPROT            => hps_h2f_lw_axi_master_arprot,        --                    .arprot
			h2f_lw_ARVALID           => hps_h2f_lw_axi_master_arvalid,       --                    .arvalid
			h2f_lw_ARREADY           => hps_h2f_lw_axi_master_arready,       --                    .arready
			h2f_lw_RID               => hps_h2f_lw_axi_master_rid,           --                    .rid
			h2f_lw_RDATA             => hps_h2f_lw_axi_master_rdata,         --                    .rdata
			h2f_lw_RRESP             => hps_h2f_lw_axi_master_rresp,         --                    .rresp
			h2f_lw_RLAST             => hps_h2f_lw_axi_master_rlast,         --                    .rlast
			h2f_lw_RVALID            => hps_h2f_lw_axi_master_rvalid,        --                    .rvalid
			h2f_lw_RREADY            => hps_h2f_lw_axi_master_rready,        --                    .rready
			f2h_irq_p0               => hps_f2h_irq0_irq,                    --            f2h_irq0.irq
			f2h_irq_p1               => hps_f2h_irq1_irq                     --            f2h_irq1.irq
		);

	jtag_uart : component soc_system_jtag_uart
		port map (
			clk            => clk_clk,                                                       --               clk.clk
			rst_n          => rst_controller_002_reset_out_reset_ports_inv,                  --             reset.reset_n
			av_chipselect  => mm_interconnect_1_jtag_uart_avalon_jtag_slave_chipselect,      -- avalon_jtag_slave.chipselect
			av_address     => mm_interconnect_1_jtag_uart_avalon_jtag_slave_address(0),      --                  .address
			av_read_n      => mm_interconnect_1_jtag_uart_avalon_jtag_slave_read_ports_inv,  --                  .read_n
			av_readdata    => mm_interconnect_1_jtag_uart_avalon_jtag_slave_readdata,        --                  .readdata
			av_write_n     => mm_interconnect_1_jtag_uart_avalon_jtag_slave_write_ports_inv, --                  .write_n
			av_writedata   => mm_interconnect_1_jtag_uart_avalon_jtag_slave_writedata,       --                  .writedata
			av_waitrequest => mm_interconnect_1_jtag_uart_avalon_jtag_slave_waitrequest,     --                  .waitrequest
			av_irq         => irq_mapper_receiver0_irq                                       --               irq.irq
		);

	master_0 : component soc_system_master_0
		generic map (
			USE_PLI     => 0,
			PLI_PORT    => 50000,
			FIFO_DEPTHS => 2
		)
		port map (
			clk_clk              => pll_using_ad1939_mclk_outclk0_clk, --          clk.clk
			clk_reset_reset      => reset_reset_n_ports_inv,           --    clk_reset.reset
			master_address       => master_0_master_address,           --       master.address
			master_readdata      => master_0_master_readdata,          --             .readdata
			master_read          => master_0_master_read,              --             .read
			master_write         => master_0_master_write,             --             .write
			master_writedata     => master_0_master_writedata,         --             .writedata
			master_waitrequest   => master_0_master_waitrequest,       --             .waitrequest
			master_readdatavalid => master_0_master_readdatavalid,     --             .readdatavalid
			master_byteenable    => master_0_master_byteenable,        --             .byteenable
			master_reset_reset   => master_0_master_reset_reset        -- master_reset.reset
		);

	onchip_memory : component soc_system_onchip_memory
		port map (
			clk        => clk_clk,                                       --   clk1.clk
			address    => mm_interconnect_0_onchip_memory_s1_address,    --     s1.address
			clken      => mm_interconnect_0_onchip_memory_s1_clken,      --       .clken
			chipselect => mm_interconnect_0_onchip_memory_s1_chipselect, --       .chipselect
			write      => mm_interconnect_0_onchip_memory_s1_write,      --       .write
			readdata   => mm_interconnect_0_onchip_memory_s1_readdata,   --       .readdata
			writedata  => mm_interconnect_0_onchip_memory_s1_writedata,  --       .writedata
			byteenable => mm_interconnect_0_onchip_memory_s1_byteenable, --       .byteenable
			reset      => rst_controller_001_reset_out_reset,            -- reset1.reset
			reset_req  => rst_controller_001_reset_out_reset_req,        --       .reset_req
			freeze     => '0'                                            -- (terminated)
		);

	pfir_testing_0 : component pFIR_Testing_dataplane_avalon
		port map (
			clk                      => pll_using_ad1939_mclk_outclk0_clk,                          --                   clock.clk
			reset                    => rst_controller_reset_out_reset,                             --                   reset.reset
			avalon_sink_valid        => avalon_st_adapter_out_0_valid,                              --   avalon_streaming_sink.valid
			avalon_sink_data         => avalon_st_adapter_out_0_data,                               --                        .data
			avalon_sink_channel      => avalon_st_adapter_out_0_channel,                            --                        .channel
			avalon_sink_error        => avalon_st_adapter_out_0_error,                              --                        .error
			avalon_source_valid      => pfir_testing_0_avalon_streaming_source_valid,               -- avalon_streaming_source.valid
			avalon_source_data       => pfir_testing_0_avalon_streaming_source_data,                --                        .data
			avalon_source_channel    => pfir_testing_0_avalon_streaming_source_channel,             --                        .channel
			avalon_source_error      => pfir_testing_0_avalon_streaming_source_error,               --                        .error
			avalon_slave_0_address   => mm_interconnect_1_pfir_testing_0_avalon_slave_0_address(0), --          avalon_slave_0.address
			avalon_slave_0_read      => mm_interconnect_1_pfir_testing_0_avalon_slave_0_read,       --                        .read
			avalon_slave_0_readdata  => mm_interconnect_1_pfir_testing_0_avalon_slave_0_readdata,   --                        .readdata
			avalon_slave_0_write     => mm_interconnect_1_pfir_testing_0_avalon_slave_0_write,      --                        .write
			avalon_slave_0_writedata => mm_interconnect_1_pfir_testing_0_avalon_slave_0_writedata,  --                        .writedata
			avalon_slave_1_address   => mm_interconnect_1_pfir_testing_0_avalon_slave_1_address,    --          avalon_slave_1.address
			avalon_slave_1_read      => mm_interconnect_1_pfir_testing_0_avalon_slave_1_read,       --                        .read
			avalon_slave_1_readdata  => mm_interconnect_1_pfir_testing_0_avalon_slave_1_readdata,   --                        .readdata
			avalon_slave_1_write     => mm_interconnect_1_pfir_testing_0_avalon_slave_1_write,      --                        .write
			avalon_slave_1_writedata => mm_interconnect_1_pfir_testing_0_avalon_slave_1_writedata   --                        .writedata
		);

	mm_interconnect_0 : component soc_system_mm_interconnect_0
		port map (
			hps_h2f_axi_master_awid                                        => hps_h2f_axi_master_awid,                       --                                       hps_h2f_axi_master.awid
			hps_h2f_axi_master_awaddr                                      => hps_h2f_axi_master_awaddr,                     --                                                         .awaddr
			hps_h2f_axi_master_awlen                                       => hps_h2f_axi_master_awlen,                      --                                                         .awlen
			hps_h2f_axi_master_awsize                                      => hps_h2f_axi_master_awsize,                     --                                                         .awsize
			hps_h2f_axi_master_awburst                                     => hps_h2f_axi_master_awburst,                    --                                                         .awburst
			hps_h2f_axi_master_awlock                                      => hps_h2f_axi_master_awlock,                     --                                                         .awlock
			hps_h2f_axi_master_awcache                                     => hps_h2f_axi_master_awcache,                    --                                                         .awcache
			hps_h2f_axi_master_awprot                                      => hps_h2f_axi_master_awprot,                     --                                                         .awprot
			hps_h2f_axi_master_awvalid                                     => hps_h2f_axi_master_awvalid,                    --                                                         .awvalid
			hps_h2f_axi_master_awready                                     => hps_h2f_axi_master_awready,                    --                                                         .awready
			hps_h2f_axi_master_wid                                         => hps_h2f_axi_master_wid,                        --                                                         .wid
			hps_h2f_axi_master_wdata                                       => hps_h2f_axi_master_wdata,                      --                                                         .wdata
			hps_h2f_axi_master_wstrb                                       => hps_h2f_axi_master_wstrb,                      --                                                         .wstrb
			hps_h2f_axi_master_wlast                                       => hps_h2f_axi_master_wlast,                      --                                                         .wlast
			hps_h2f_axi_master_wvalid                                      => hps_h2f_axi_master_wvalid,                     --                                                         .wvalid
			hps_h2f_axi_master_wready                                      => hps_h2f_axi_master_wready,                     --                                                         .wready
			hps_h2f_axi_master_bid                                         => hps_h2f_axi_master_bid,                        --                                                         .bid
			hps_h2f_axi_master_bresp                                       => hps_h2f_axi_master_bresp,                      --                                                         .bresp
			hps_h2f_axi_master_bvalid                                      => hps_h2f_axi_master_bvalid,                     --                                                         .bvalid
			hps_h2f_axi_master_bready                                      => hps_h2f_axi_master_bready,                     --                                                         .bready
			hps_h2f_axi_master_arid                                        => hps_h2f_axi_master_arid,                       --                                                         .arid
			hps_h2f_axi_master_araddr                                      => hps_h2f_axi_master_araddr,                     --                                                         .araddr
			hps_h2f_axi_master_arlen                                       => hps_h2f_axi_master_arlen,                      --                                                         .arlen
			hps_h2f_axi_master_arsize                                      => hps_h2f_axi_master_arsize,                     --                                                         .arsize
			hps_h2f_axi_master_arburst                                     => hps_h2f_axi_master_arburst,                    --                                                         .arburst
			hps_h2f_axi_master_arlock                                      => hps_h2f_axi_master_arlock,                     --                                                         .arlock
			hps_h2f_axi_master_arcache                                     => hps_h2f_axi_master_arcache,                    --                                                         .arcache
			hps_h2f_axi_master_arprot                                      => hps_h2f_axi_master_arprot,                     --                                                         .arprot
			hps_h2f_axi_master_arvalid                                     => hps_h2f_axi_master_arvalid,                    --                                                         .arvalid
			hps_h2f_axi_master_arready                                     => hps_h2f_axi_master_arready,                    --                                                         .arready
			hps_h2f_axi_master_rid                                         => hps_h2f_axi_master_rid,                        --                                                         .rid
			hps_h2f_axi_master_rdata                                       => hps_h2f_axi_master_rdata,                      --                                                         .rdata
			hps_h2f_axi_master_rresp                                       => hps_h2f_axi_master_rresp,                      --                                                         .rresp
			hps_h2f_axi_master_rlast                                       => hps_h2f_axi_master_rlast,                      --                                                         .rlast
			hps_h2f_axi_master_rvalid                                      => hps_h2f_axi_master_rvalid,                     --                                                         .rvalid
			hps_h2f_axi_master_rready                                      => hps_h2f_axi_master_rready,                     --                                                         .rready
			clk_hps_clk_clk                                                => clk_clk,                                       --                                              clk_hps_clk.clk
			hps_h2f_axi_master_agent_clk_reset_reset_bridge_in_reset_reset => rst_controller_003_reset_out_reset,            -- hps_h2f_axi_master_agent_clk_reset_reset_bridge_in_reset.reset
			onchip_memory_reset1_reset_bridge_in_reset_reset               => rst_controller_001_reset_out_reset,            --               onchip_memory_reset1_reset_bridge_in_reset.reset
			onchip_memory_s1_address                                       => mm_interconnect_0_onchip_memory_s1_address,    --                                         onchip_memory_s1.address
			onchip_memory_s1_write                                         => mm_interconnect_0_onchip_memory_s1_write,      --                                                         .write
			onchip_memory_s1_readdata                                      => mm_interconnect_0_onchip_memory_s1_readdata,   --                                                         .readdata
			onchip_memory_s1_writedata                                     => mm_interconnect_0_onchip_memory_s1_writedata,  --                                                         .writedata
			onchip_memory_s1_byteenable                                    => mm_interconnect_0_onchip_memory_s1_byteenable, --                                                         .byteenable
			onchip_memory_s1_chipselect                                    => mm_interconnect_0_onchip_memory_s1_chipselect, --                                                         .chipselect
			onchip_memory_s1_clken                                         => mm_interconnect_0_onchip_memory_s1_clken       --                                                         .clken
		);

	mm_interconnect_1 : component soc_system_mm_interconnect_1
		port map (
			hps_h2f_lw_axi_master_awid                                        => hps_h2f_lw_axi_master_awid,                                --                                       hps_h2f_lw_axi_master.awid
			hps_h2f_lw_axi_master_awaddr                                      => hps_h2f_lw_axi_master_awaddr,                              --                                                            .awaddr
			hps_h2f_lw_axi_master_awlen                                       => hps_h2f_lw_axi_master_awlen,                               --                                                            .awlen
			hps_h2f_lw_axi_master_awsize                                      => hps_h2f_lw_axi_master_awsize,                              --                                                            .awsize
			hps_h2f_lw_axi_master_awburst                                     => hps_h2f_lw_axi_master_awburst,                             --                                                            .awburst
			hps_h2f_lw_axi_master_awlock                                      => hps_h2f_lw_axi_master_awlock,                              --                                                            .awlock
			hps_h2f_lw_axi_master_awcache                                     => hps_h2f_lw_axi_master_awcache,                             --                                                            .awcache
			hps_h2f_lw_axi_master_awprot                                      => hps_h2f_lw_axi_master_awprot,                              --                                                            .awprot
			hps_h2f_lw_axi_master_awvalid                                     => hps_h2f_lw_axi_master_awvalid,                             --                                                            .awvalid
			hps_h2f_lw_axi_master_awready                                     => hps_h2f_lw_axi_master_awready,                             --                                                            .awready
			hps_h2f_lw_axi_master_wid                                         => hps_h2f_lw_axi_master_wid,                                 --                                                            .wid
			hps_h2f_lw_axi_master_wdata                                       => hps_h2f_lw_axi_master_wdata,                               --                                                            .wdata
			hps_h2f_lw_axi_master_wstrb                                       => hps_h2f_lw_axi_master_wstrb,                               --                                                            .wstrb
			hps_h2f_lw_axi_master_wlast                                       => hps_h2f_lw_axi_master_wlast,                               --                                                            .wlast
			hps_h2f_lw_axi_master_wvalid                                      => hps_h2f_lw_axi_master_wvalid,                              --                                                            .wvalid
			hps_h2f_lw_axi_master_wready                                      => hps_h2f_lw_axi_master_wready,                              --                                                            .wready
			hps_h2f_lw_axi_master_bid                                         => hps_h2f_lw_axi_master_bid,                                 --                                                            .bid
			hps_h2f_lw_axi_master_bresp                                       => hps_h2f_lw_axi_master_bresp,                               --                                                            .bresp
			hps_h2f_lw_axi_master_bvalid                                      => hps_h2f_lw_axi_master_bvalid,                              --                                                            .bvalid
			hps_h2f_lw_axi_master_bready                                      => hps_h2f_lw_axi_master_bready,                              --                                                            .bready
			hps_h2f_lw_axi_master_arid                                        => hps_h2f_lw_axi_master_arid,                                --                                                            .arid
			hps_h2f_lw_axi_master_araddr                                      => hps_h2f_lw_axi_master_araddr,                              --                                                            .araddr
			hps_h2f_lw_axi_master_arlen                                       => hps_h2f_lw_axi_master_arlen,                               --                                                            .arlen
			hps_h2f_lw_axi_master_arsize                                      => hps_h2f_lw_axi_master_arsize,                              --                                                            .arsize
			hps_h2f_lw_axi_master_arburst                                     => hps_h2f_lw_axi_master_arburst,                             --                                                            .arburst
			hps_h2f_lw_axi_master_arlock                                      => hps_h2f_lw_axi_master_arlock,                              --                                                            .arlock
			hps_h2f_lw_axi_master_arcache                                     => hps_h2f_lw_axi_master_arcache,                             --                                                            .arcache
			hps_h2f_lw_axi_master_arprot                                      => hps_h2f_lw_axi_master_arprot,                              --                                                            .arprot
			hps_h2f_lw_axi_master_arvalid                                     => hps_h2f_lw_axi_master_arvalid,                             --                                                            .arvalid
			hps_h2f_lw_axi_master_arready                                     => hps_h2f_lw_axi_master_arready,                             --                                                            .arready
			hps_h2f_lw_axi_master_rid                                         => hps_h2f_lw_axi_master_rid,                                 --                                                            .rid
			hps_h2f_lw_axi_master_rdata                                       => hps_h2f_lw_axi_master_rdata,                               --                                                            .rdata
			hps_h2f_lw_axi_master_rresp                                       => hps_h2f_lw_axi_master_rresp,                               --                                                            .rresp
			hps_h2f_lw_axi_master_rlast                                       => hps_h2f_lw_axi_master_rlast,                               --                                                            .rlast
			hps_h2f_lw_axi_master_rvalid                                      => hps_h2f_lw_axi_master_rvalid,                              --                                                            .rvalid
			hps_h2f_lw_axi_master_rready                                      => hps_h2f_lw_axi_master_rready,                              --                                                            .rready
			clk_hps_clk_clk                                                   => clk_clk,                                                   --                                                 clk_hps_clk.clk
			PLL_using_AD1939_MCLK_outclk0_clk                                 => pll_using_ad1939_mclk_outclk0_clk,                         --                               PLL_using_AD1939_MCLK_outclk0.clk
			hps_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset_reset => rst_controller_003_reset_out_reset,                        -- hps_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset.reset
			jtag_uart_reset_reset_bridge_in_reset_reset                       => rst_controller_002_reset_out_reset,                        --                       jtag_uart_reset_reset_bridge_in_reset.reset
			master_0_clk_reset_reset_bridge_in_reset_reset                    => rst_controller_reset_out_reset,                            --                    master_0_clk_reset_reset_bridge_in_reset.reset
			pFIR_Testing_0_reset_reset_bridge_in_reset_reset                  => rst_controller_reset_out_reset,                            --                  pFIR_Testing_0_reset_reset_bridge_in_reset.reset
			SystemID_reset_reset_bridge_in_reset_reset                        => rst_controller_001_reset_out_reset,                        --                        SystemID_reset_reset_bridge_in_reset.reset
			master_0_master_address                                           => master_0_master_address,                                   --                                             master_0_master.address
			master_0_master_waitrequest                                       => master_0_master_waitrequest,                               --                                                            .waitrequest
			master_0_master_byteenable                                        => master_0_master_byteenable,                                --                                                            .byteenable
			master_0_master_read                                              => master_0_master_read,                                      --                                                            .read
			master_0_master_readdata                                          => master_0_master_readdata,                                  --                                                            .readdata
			master_0_master_readdatavalid                                     => master_0_master_readdatavalid,                             --                                                            .readdatavalid
			master_0_master_write                                             => master_0_master_write,                                     --                                                            .write
			master_0_master_writedata                                         => master_0_master_writedata,                                 --                                                            .writedata
			jtag_uart_avalon_jtag_slave_address                               => mm_interconnect_1_jtag_uart_avalon_jtag_slave_address,     --                                 jtag_uart_avalon_jtag_slave.address
			jtag_uart_avalon_jtag_slave_write                                 => mm_interconnect_1_jtag_uart_avalon_jtag_slave_write,       --                                                            .write
			jtag_uart_avalon_jtag_slave_read                                  => mm_interconnect_1_jtag_uart_avalon_jtag_slave_read,        --                                                            .read
			jtag_uart_avalon_jtag_slave_readdata                              => mm_interconnect_1_jtag_uart_avalon_jtag_slave_readdata,    --                                                            .readdata
			jtag_uart_avalon_jtag_slave_writedata                             => mm_interconnect_1_jtag_uart_avalon_jtag_slave_writedata,   --                                                            .writedata
			jtag_uart_avalon_jtag_slave_waitrequest                           => mm_interconnect_1_jtag_uart_avalon_jtag_slave_waitrequest, --                                                            .waitrequest
			jtag_uart_avalon_jtag_slave_chipselect                            => mm_interconnect_1_jtag_uart_avalon_jtag_slave_chipselect,  --                                                            .chipselect
			pFIR_Testing_0_avalon_slave_0_address                             => mm_interconnect_1_pfir_testing_0_avalon_slave_0_address,   --                               pFIR_Testing_0_avalon_slave_0.address
			pFIR_Testing_0_avalon_slave_0_write                               => mm_interconnect_1_pfir_testing_0_avalon_slave_0_write,     --                                                            .write
			pFIR_Testing_0_avalon_slave_0_read                                => mm_interconnect_1_pfir_testing_0_avalon_slave_0_read,      --                                                            .read
			pFIR_Testing_0_avalon_slave_0_readdata                            => mm_interconnect_1_pfir_testing_0_avalon_slave_0_readdata,  --                                                            .readdata
			pFIR_Testing_0_avalon_slave_0_writedata                           => mm_interconnect_1_pfir_testing_0_avalon_slave_0_writedata, --                                                            .writedata
			pFIR_Testing_0_avalon_slave_1_address                             => mm_interconnect_1_pfir_testing_0_avalon_slave_1_address,   --                               pFIR_Testing_0_avalon_slave_1.address
			pFIR_Testing_0_avalon_slave_1_write                               => mm_interconnect_1_pfir_testing_0_avalon_slave_1_write,     --                                                            .write
			pFIR_Testing_0_avalon_slave_1_read                                => mm_interconnect_1_pfir_testing_0_avalon_slave_1_read,      --                                                            .read
			pFIR_Testing_0_avalon_slave_1_readdata                            => mm_interconnect_1_pfir_testing_0_avalon_slave_1_readdata,  --                                                            .readdata
			pFIR_Testing_0_avalon_slave_1_writedata                           => mm_interconnect_1_pfir_testing_0_avalon_slave_1_writedata, --                                                            .writedata
			SystemID_control_slave_address                                    => mm_interconnect_1_systemid_control_slave_address,          --                                      SystemID_control_slave.address
			SystemID_control_slave_readdata                                   => mm_interconnect_1_systemid_control_slave_readdata          --                                                            .readdata
		);

	irq_mapper : component soc_system_irq_mapper
		port map (
			clk           => open,                     --       clk.clk
			reset         => open,                     -- clk_reset.reset
			receiver0_irq => irq_mapper_receiver0_irq, -- receiver0.irq
			sender_irq    => hps_f2h_irq0_irq          --    sender.irq
		);

	irq_mapper_001 : component soc_system_irq_mapper_001
		port map (
			clk        => open,             --       clk.clk
			reset      => open,             -- clk_reset.reset
			sender_irq => hps_f2h_irq1_irq  --    sender.irq
		);

	avalon_st_adapter : component soc_system_avalon_st_adapter
		generic map (
			inBitsPerSymbol => 32,
			inUsePackets    => 0,
			inDataWidth     => 32,
			inChannelWidth  => 2,
			inErrorWidth    => 2,
			inUseEmptyPort  => 0,
			inUseValid      => 1,
			inUseReady      => 0,
			inReadyLatency  => 0,
			outDataWidth    => 32,
			outChannelWidth => 2,
			outErrorWidth   => 2,
			outUseEmptyPort => 0,
			outUseValid     => 1,
			outUseReady     => 0,
			outReadyLatency => 0
		)
		port map (
			in_clk_0_clk   => pll_using_ad1939_mclk_outclk0_clk,              -- in_clk_0.clk
			in_rst_0_reset => rst_controller_reset_out_reset,                 -- in_rst_0.reset
			in_0_data      => fe_qsys_ad1939_audio_mini_v1_0_line_in_data,    --     in_0.data
			in_0_valid     => fe_qsys_ad1939_audio_mini_v1_0_line_in_valid,   --         .valid
			in_0_error     => fe_qsys_ad1939_audio_mini_v1_0_line_in_error,   --         .error
			in_0_channel   => fe_qsys_ad1939_audio_mini_v1_0_line_in_channel, --         .channel
			out_0_data     => avalon_st_adapter_out_0_data,                   --    out_0.data
			out_0_valid    => avalon_st_adapter_out_0_valid,                  --         .valid
			out_0_error    => avalon_st_adapter_out_0_error,                  --         .error
			out_0_channel  => avalon_st_adapter_out_0_channel                 --         .channel
		);

	avalon_st_adapter_001 : component soc_system_avalon_st_adapter_001
		generic map (
			inBitsPerSymbol => 32,
			inUsePackets    => 0,
			inDataWidth     => 32,
			inChannelWidth  => 2,
			inErrorWidth    => 2,
			inUseEmptyPort  => 0,
			inUseValid      => 1,
			inUseReady      => 0,
			inReadyLatency  => 0,
			outDataWidth    => 32,
			outChannelWidth => 2,
			outErrorWidth   => 2,
			outUseEmptyPort => 0,
			outUseValid     => 1,
			outUseReady     => 0,
			outReadyLatency => 0
		)
		port map (
			in_clk_0_clk   => pll_using_ad1939_mclk_outclk0_clk,              -- in_clk_0.clk
			in_rst_0_reset => rst_controller_reset_out_reset,                 -- in_rst_0.reset
			in_0_data      => pfir_testing_0_avalon_streaming_source_data,    --     in_0.data
			in_0_valid     => pfir_testing_0_avalon_streaming_source_valid,   --         .valid
			in_0_error     => pfir_testing_0_avalon_streaming_source_error,   --         .error
			in_0_channel   => pfir_testing_0_avalon_streaming_source_channel, --         .channel
			out_0_data     => avalon_st_adapter_001_out_0_data,               --    out_0.data
			out_0_valid    => avalon_st_adapter_001_out_0_valid,              --         .valid
			out_0_error    => avalon_st_adapter_001_out_0_error,              --         .error
			out_0_channel  => avalon_st_adapter_001_out_0_channel             --         .channel
		);

	rst_controller : component soc_system_rst_controller
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,           -- reset_in0.reset
			clk            => pll_using_ad1939_mclk_outclk0_clk, --       clk.clk
			reset_out      => rst_controller_reset_out_reset,    -- reset_out.reset
			reset_req      => open,                              -- (terminated)
			reset_req_in0  => '0',                               -- (terminated)
			reset_in1      => '0',                               -- (terminated)
			reset_req_in1  => '0',                               -- (terminated)
			reset_in2      => '0',                               -- (terminated)
			reset_req_in2  => '0',                               -- (terminated)
			reset_in3      => '0',                               -- (terminated)
			reset_req_in3  => '0',                               -- (terminated)
			reset_in4      => '0',                               -- (terminated)
			reset_req_in4  => '0',                               -- (terminated)
			reset_in5      => '0',                               -- (terminated)
			reset_req_in5  => '0',                               -- (terminated)
			reset_in6      => '0',                               -- (terminated)
			reset_req_in6  => '0',                               -- (terminated)
			reset_in7      => '0',                               -- (terminated)
			reset_req_in7  => '0',                               -- (terminated)
			reset_in8      => '0',                               -- (terminated)
			reset_req_in8  => '0',                               -- (terminated)
			reset_in9      => '0',                               -- (terminated)
			reset_req_in9  => '0',                               -- (terminated)
			reset_in10     => '0',                               -- (terminated)
			reset_req_in10 => '0',                               -- (terminated)
			reset_in11     => '0',                               -- (terminated)
			reset_req_in11 => '0',                               -- (terminated)
			reset_in12     => '0',                               -- (terminated)
			reset_req_in12 => '0',                               -- (terminated)
			reset_in13     => '0',                               -- (terminated)
			reset_req_in13 => '0',                               -- (terminated)
			reset_in14     => '0',                               -- (terminated)
			reset_req_in14 => '0',                               -- (terminated)
			reset_in15     => '0',                               -- (terminated)
			reset_req_in15 => '0'                                -- (terminated)
		);

	rst_controller_001 : component soc_system_rst_controller_001
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 1,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,                -- reset_in0.reset
			clk            => clk_clk,                                --       clk.clk
			reset_out      => rst_controller_001_reset_out_reset,     -- reset_out.reset
			reset_req      => rst_controller_001_reset_out_reset_req, --          .reset_req
			reset_req_in0  => '0',                                    -- (terminated)
			reset_in1      => '0',                                    -- (terminated)
			reset_req_in1  => '0',                                    -- (terminated)
			reset_in2      => '0',                                    -- (terminated)
			reset_req_in2  => '0',                                    -- (terminated)
			reset_in3      => '0',                                    -- (terminated)
			reset_req_in3  => '0',                                    -- (terminated)
			reset_in4      => '0',                                    -- (terminated)
			reset_req_in4  => '0',                                    -- (terminated)
			reset_in5      => '0',                                    -- (terminated)
			reset_req_in5  => '0',                                    -- (terminated)
			reset_in6      => '0',                                    -- (terminated)
			reset_req_in6  => '0',                                    -- (terminated)
			reset_in7      => '0',                                    -- (terminated)
			reset_req_in7  => '0',                                    -- (terminated)
			reset_in8      => '0',                                    -- (terminated)
			reset_req_in8  => '0',                                    -- (terminated)
			reset_in9      => '0',                                    -- (terminated)
			reset_req_in9  => '0',                                    -- (terminated)
			reset_in10     => '0',                                    -- (terminated)
			reset_req_in10 => '0',                                    -- (terminated)
			reset_in11     => '0',                                    -- (terminated)
			reset_req_in11 => '0',                                    -- (terminated)
			reset_in12     => '0',                                    -- (terminated)
			reset_req_in12 => '0',                                    -- (terminated)
			reset_in13     => '0',                                    -- (terminated)
			reset_req_in13 => '0',                                    -- (terminated)
			reset_in14     => '0',                                    -- (terminated)
			reset_req_in14 => '0',                                    -- (terminated)
			reset_in15     => '0',                                    -- (terminated)
			reset_req_in15 => '0'                                     -- (terminated)
		);

	rst_controller_002 : component soc_system_rst_controller_002
		generic map (
			NUM_RESET_INPUTS          => 2,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,            -- reset_in0.reset
			reset_in1      => master_0_master_reset_reset,        -- reset_in1.reset
			clk            => clk_clk,                            --       clk.clk
			reset_out      => rst_controller_002_reset_out_reset, -- reset_out.reset
			reset_req      => open,                               -- (terminated)
			reset_req_in0  => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_in2      => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	rst_controller_003 : component soc_system_rst_controller
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => hps_h2f_reset_reset_n_ports_inv,    -- reset_in0.reset
			clk            => clk_clk,                            --       clk.clk
			reset_out      => rst_controller_003_reset_out_reset, -- reset_out.reset
			reset_req      => open,                               -- (terminated)
			reset_req_in0  => '0',                                -- (terminated)
			reset_in1      => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_in2      => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	hps_h2f_reset_reset_n_ports_inv <= not hps_h2f_reset_reset;

	reset_reset_n_ports_inv <= not reset_reset_n;

	mm_interconnect_1_jtag_uart_avalon_jtag_slave_read_ports_inv <= not mm_interconnect_1_jtag_uart_avalon_jtag_slave_read;

	mm_interconnect_1_jtag_uart_avalon_jtag_slave_write_ports_inv <= not mm_interconnect_1_jtag_uart_avalon_jtag_slave_write;

	rst_controller_001_reset_out_reset_ports_inv <= not rst_controller_001_reset_out_reset;

	rst_controller_002_reset_out_reset_ports_inv <= not rst_controller_002_reset_out_reset;

	hps_h2f_reset_reset_n <= hps_h2f_reset_reset;

end architecture rtl; -- of soc_system
