-- pll_sys.vhd

-- Generated using ACDS version 18.0 614

library IEEE;
library pll_sys_altera_iopll_180;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity pll_sys is
	port (
		locked   : out std_logic;        --  locked.export
		outclk_0 : out std_logic;        -- outclk0.clk
		refclk   : in  std_logic := '0'; --  refclk.clk
		rst      : in  std_logic := '0'  --   reset.reset
	);
end entity pll_sys;

architecture rtl of pll_sys is
	component pll_sys_altera_iopll_180_hm2x5zi is
		port (
			rst      : in  std_logic := 'X'; -- reset
			refclk   : in  std_logic := 'X'; -- clk
			locked   : out std_logic;        -- export
			outclk_0 : out std_logic         -- clk
		);
	end component pll_sys_altera_iopll_180_hm2x5zi;

	for iopll_0 : pll_sys_altera_iopll_180_hm2x5zi
		use entity pll_sys_altera_iopll_180.pll_sys_altera_iopll_180_hm2x5zi;
begin

	iopll_0 : component pll_sys_altera_iopll_180_hm2x5zi
		port map (
			rst      => rst,      --   reset.reset
			refclk   => refclk,   --  refclk.clk
			locked   => locked,   --  locked.export
			outclk_0 => outclk_0  -- outclk0.clk
		);

end architecture rtl; -- of pll_sys
