----------------------------------------------------------------------------------------------------
-- Copyright (c) ReFLEX CES 1998-2016
--
-- Use of this source code through a simulator and/or a compiler tool
-- is illegal if not authorised through ReFLEX CES License agreement.
----------------------------------------------------------------------------------------------------
----------------------------------------------------------------------------------------------------
-- Author      : Fr�d�ric Lavenant       flavenant@reflexces.com
-- Company     : ReFLEX CES
--               2, rue du gevaudan
--               91047 LISSES
--               FRANCE
--               http://www.reflexces.com
----------------------------------------------------------------------------------------------------
-- Description :
-- Duplicate input to outputs.
-- Input is ready only if all outputs are ready. 
--
----------------------------------------------------------------------------------------------------
-- Version      Date            Author               Description
-- 0.1          2014/01/28      FLA                  Creation
-- 0.2          2016/10/13      JDU                 Change lib_jlf to work 
----------------------------------------------------------------------------------------------------
library ieee;
use     ieee.std_logic_1164.all;
use     ieee.numeric_std.all;

library work;
use     work.pkg_std.all;
use     work.pkg_std_unsigned.all;

entity bus_duplicate is
    generic (
          NB_OUTPUT         : integer           := 4                        -- Number of inputs to manage
        ; DATA_WIDTH        : integer           := 33                       -- Input is NB_OUTPUT*DATA_WIDTH
    );              
    port (              
          rst               : in    sl                                      -- Active high (A)synchronous reset
        ; clk               : in    sl                                      -- Clock
            
        ; i_dat             : in    slv(DATA_WIDTH-1 downto 0)              -- Input data 
        ; i_vld             : in    sl                                      -- Valid input
        ; i_rdy             : out   sl                                      -- Input ready
            
        ; o_dat             : out   slv(NB_OUTPUT*DATA_WIDTH-1 downto 0)    -- Output data
        ; o_vld             : out   slv(NB_OUTPUT-1 downto 0)               -- Output valid
        ; o_rdy             : in    slv(NB_OUTPUT-1 downto 0)               -- Output ready
    );
end entity bus_duplicate;

architecture rtl of bus_duplicate is
    --============================================================================================================================
    -- Function and Procedure declarations
    --============================================================================================================================
    
    --============================================================================================================================
    -- Constant and Type declarations
    --============================================================================================================================

    --============================================================================================================================
    -- Component declarations
    --============================================================================================================================
    
    --============================================================================================================================
    -- Signal declarations
    --============================================================================================================================
    signal s_o_dat  : slv(DATA_WIDTH-1 downto 0);
    signal s_o_vld  : slv(NB_OUTPUT-1 downto 0);
    signal s_i_rdy  : sl;
begin
    --############################################################################################################################
    --############################################################################################################################
    -- Generate output
    --############################################################################################################################
    --############################################################################################################################
    --============================================================================================================================
    -- Process
    --============================================================================================================================
    gen_output : for i in 0 to NB_OUTPUT-1 generate
    begin
        ------------------------------------------------
        -- For valid
        ------------------------------------------------
        process (rst, clk)
        begin
        if rst='1' then
            s_o_vld(i) <= '0';
        elsif rising_edge(clk) then
            if (s_o_vld(i)='0' or o_rdy(i)='1') then s_o_vld(i) <= i_vld and s_i_rdy; end if;
        end if;
        end process;
        
        ------------------------------------------------
        -- For data
        ------------------------------------------------
        o_dat((i+1)*DATA_WIDTH-1 downto i*DATA_WIDTH) <= s_o_dat;
    end generate gen_output;
    
    --============================================================================================================================
    -- Assignment
    --============================================================================================================================
    o_vld <= s_o_vld;
    
    --############################################################################################################################
    --############################################################################################################################
    -- Generate output data
    --############################################################################################################################
    --############################################################################################################################
    process (rst, clk)
    begin
    if rst='1' then
        s_o_dat   <= (others=>'0');
    elsif rising_edge(clk) then
        if i_vld='1' and s_i_rdy='1' then s_o_dat <= i_dat; end if;
    end if;
    end process;
    
    --############################################################################################################################
    --############################################################################################################################
    -- Generate input ready 
    --############################################################################################################################
    --############################################################################################################################
    s_i_rdy <= '1' when or1(s_o_vld)='0'    else    -- all outputs are not valid
               '1' when and1(o_rdy)='1'     else    -- all outputs are ready
               '0';
    i_rdy   <= s_i_rdy;
end architecture rtl;
