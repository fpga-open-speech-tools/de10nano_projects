AD1939_reg_init_ROM_inst : AD1939_reg_init_ROM PORT MAP (
		address	 => address_sig,
		clock	 => clock_sig,
		q	 => q_sig
	);
