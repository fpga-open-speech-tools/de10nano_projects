/*--------------------------------------------------------------------------------------------------------------------------------------------------------------
Author      : Jean-Louis FLOQUET
Title       : Package for usual constants
File        : pkg_cst.vhd
Application : RTL & Simulation
Created     : 2007, June 5th
Last update : 2013/12/19 14:55
Version     : 1.05.01
Dependency  : pkg_std
----------------------------------------------------------------------------------------------------------------------------------------------------------------
Description : This package contains usefull constants
----------------------------------------------------------------------------------------------------------------------------------------------------------------
   Rev.  |    Date    | Description
 1.05.01 | 2013/12/19 | 1) Chg : VHDL-2008 required
 1.04.01 | 2013/06/17 | 1) New : Add XS_xx up to 1024
 1.03.01 | 2011/10/25 | 1) New : Add ZEROS_xx and ONES_xx up to 1024
 1.02.01 | 2011/09/30 | 1) New : Add ZEROS_xx and ONES_xx up to 256
 1.01.01 | 2007/08/30 | 1) New : Some mathematical constants
 1.00.00 | 2007/06/05 | Initial Release
         |            |
--------------------------------------------------------------------------------------------------------------------------------------------------------------*/
library ieee;
use     ieee.std_logic_1164.all;
use     ieee.numeric_std.all;

library work;
use     work.pkg_std.all;

package pkg_cst is
--**************************************************************************************************************************************************************
-- ZERO
--**************************************************************************************************************************************************************
	constant ZEROS      : slv(1023 downto 0) := (others=>'0');
	constant ZEROS_1    : slv1    := (others=>'0'); constant ZEROS_2    : slv2    := (others=>'0'); constant ZEROS_3    : slv3    := (others=>'0'); constant ZEROS_4    : slv4    := (others=>'0');
	constant ZEROS_5    : slv5    := (others=>'0'); constant ZEROS_6    : slv6    := (others=>'0'); constant ZEROS_7    : slv7    := (others=>'0'); constant ZEROS_8    : slv8    := (others=>'0');
	constant ZEROS_9    : slv9    := (others=>'0'); constant ZEROS_10   : slv10   := (others=>'0'); constant ZEROS_11   : slv11   := (others=>'0'); constant ZEROS_12   : slv12   := (others=>'0');
	constant ZEROS_13   : slv13   := (others=>'0'); constant ZEROS_14   : slv14   := (others=>'0'); constant ZEROS_15   : slv15   := (others=>'0'); constant ZEROS_16   : slv16   := (others=>'0');
	constant ZEROS_17   : slv17   := (others=>'0'); constant ZEROS_18   : slv18   := (others=>'0'); constant ZEROS_19   : slv19   := (others=>'0'); constant ZEROS_20   : slv20   := (others=>'0');
	constant ZEROS_21   : slv21   := (others=>'0'); constant ZEROS_22   : slv22   := (others=>'0'); constant ZEROS_23   : slv23   := (others=>'0'); constant ZEROS_24   : slv24   := (others=>'0');
	constant ZEROS_25   : slv25   := (others=>'0'); constant ZEROS_26   : slv26   := (others=>'0'); constant ZEROS_27   : slv27   := (others=>'0'); constant ZEROS_28   : slv28   := (others=>'0');
	constant ZEROS_29   : slv29   := (others=>'0'); constant ZEROS_30   : slv30   := (others=>'0'); constant ZEROS_31   : slv31   := (others=>'0'); constant ZEROS_32   : slv32   := (others=>'0');
	constant ZEROS_33   : slv33   := (others=>'0'); constant ZEROS_34   : slv34   := (others=>'0'); constant ZEROS_35   : slv35   := (others=>'0'); constant ZEROS_36   : slv36   := (others=>'0');
	constant ZEROS_37   : slv37   := (others=>'0'); constant ZEROS_38   : slv38   := (others=>'0'); constant ZEROS_39   : slv39   := (others=>'0'); constant ZEROS_40   : slv40   := (others=>'0');
	constant ZEROS_41   : slv41   := (others=>'0'); constant ZEROS_42   : slv42   := (others=>'0'); constant ZEROS_43   : slv43   := (others=>'0'); constant ZEROS_44   : slv44   := (others=>'0');
	constant ZEROS_45   : slv45   := (others=>'0'); constant ZEROS_46   : slv46   := (others=>'0'); constant ZEROS_47   : slv47   := (others=>'0'); constant ZEROS_48   : slv48   := (others=>'0');
	constant ZEROS_49   : slv49   := (others=>'0'); constant ZEROS_50   : slv50   := (others=>'0'); constant ZEROS_51   : slv51   := (others=>'0'); constant ZEROS_52   : slv52   := (others=>'0');
	constant ZEROS_53   : slv53   := (others=>'0'); constant ZEROS_54   : slv54   := (others=>'0'); constant ZEROS_55   : slv55   := (others=>'0'); constant ZEROS_56   : slv56   := (others=>'0');
	constant ZEROS_57   : slv57   := (others=>'0'); constant ZEROS_58   : slv58   := (others=>'0'); constant ZEROS_59   : slv59   := (others=>'0'); constant ZEROS_60   : slv60   := (others=>'0');
	constant ZEROS_61   : slv61   := (others=>'0'); constant ZEROS_62   : slv62   := (others=>'0'); constant ZEROS_63   : slv63   := (others=>'0'); constant ZEROS_64   : slv64   := (others=>'0');
	constant ZEROS_65   : slv65   := (others=>'0'); constant ZEROS_66   : slv66   := (others=>'0'); constant ZEROS_67   : slv67   := (others=>'0'); constant ZEROS_68   : slv68   := (others=>'0');
	constant ZEROS_69   : slv69   := (others=>'0'); constant ZEROS_70   : slv70   := (others=>'0'); constant ZEROS_71   : slv71   := (others=>'0'); constant ZEROS_72   : slv72   := (others=>'0');
	constant ZEROS_73   : slv73   := (others=>'0'); constant ZEROS_74   : slv74   := (others=>'0'); constant ZEROS_75   : slv75   := (others=>'0'); constant ZEROS_76   : slv76   := (others=>'0');
	constant ZEROS_77   : slv77   := (others=>'0'); constant ZEROS_78   : slv78   := (others=>'0'); constant ZEROS_79   : slv79   := (others=>'0'); constant ZEROS_80   : slv80   := (others=>'0');
	constant ZEROS_81   : slv81   := (others=>'0'); constant ZEROS_82   : slv82   := (others=>'0'); constant ZEROS_83   : slv83   := (others=>'0'); constant ZEROS_84   : slv84   := (others=>'0');
	constant ZEROS_85   : slv85   := (others=>'0'); constant ZEROS_86   : slv86   := (others=>'0'); constant ZEROS_87   : slv87   := (others=>'0'); constant ZEROS_88   : slv88   := (others=>'0');
	constant ZEROS_89   : slv89   := (others=>'0'); constant ZEROS_90   : slv90   := (others=>'0'); constant ZEROS_91   : slv91   := (others=>'0'); constant ZEROS_92   : slv92   := (others=>'0');
	constant ZEROS_93   : slv93   := (others=>'0'); constant ZEROS_94   : slv94   := (others=>'0'); constant ZEROS_95   : slv95   := (others=>'0'); constant ZEROS_96   : slv96   := (others=>'0');
	constant ZEROS_97   : slv97   := (others=>'0'); constant ZEROS_98   : slv98   := (others=>'0'); constant ZEROS_99   : slv99   := (others=>'0'); constant ZEROS_100  : slv100  := (others=>'0');
	constant ZEROS_101  : slv101  := (others=>'0'); constant ZEROS_102  : slv102  := (others=>'0'); constant ZEROS_103  : slv103  := (others=>'0'); constant ZEROS_104  : slv104  := (others=>'0');
	constant ZEROS_105  : slv105  := (others=>'0'); constant ZEROS_106  : slv106  := (others=>'0'); constant ZEROS_107  : slv107  := (others=>'0'); constant ZEROS_108  : slv108  := (others=>'0');
	constant ZEROS_109  : slv109  := (others=>'0'); constant ZEROS_110  : slv110  := (others=>'0'); constant ZEROS_111  : slv111  := (others=>'0'); constant ZEROS_112  : slv112  := (others=>'0');
	constant ZEROS_113  : slv113  := (others=>'0'); constant ZEROS_114  : slv114  := (others=>'0'); constant ZEROS_115  : slv115  := (others=>'0'); constant ZEROS_116  : slv116  := (others=>'0');
	constant ZEROS_117  : slv117  := (others=>'0'); constant ZEROS_118  : slv118  := (others=>'0'); constant ZEROS_119  : slv119  := (others=>'0'); constant ZEROS_120  : slv120  := (others=>'0');
	constant ZEROS_121  : slv121  := (others=>'0'); constant ZEROS_122  : slv122  := (others=>'0'); constant ZEROS_123  : slv123  := (others=>'0'); constant ZEROS_124  : slv124  := (others=>'0');
	constant ZEROS_125  : slv125  := (others=>'0'); constant ZEROS_126  : slv126  := (others=>'0'); constant ZEROS_127  : slv127  := (others=>'0'); constant ZEROS_128  : slv128  := (others=>'0');
	constant ZEROS_129  : slv129  := (others=>'0'); constant ZEROS_130  : slv130  := (others=>'0'); constant ZEROS_131  : slv131  := (others=>'0'); constant ZEROS_132  : slv132  := (others=>'0');
	constant ZEROS_133  : slv133  := (others=>'0'); constant ZEROS_134  : slv134  := (others=>'0'); constant ZEROS_135  : slv135  := (others=>'0'); constant ZEROS_136  : slv136  := (others=>'0');
	constant ZEROS_137  : slv137  := (others=>'0'); constant ZEROS_138  : slv138  := (others=>'0'); constant ZEROS_139  : slv139  := (others=>'0'); constant ZEROS_140  : slv140  := (others=>'0');
	constant ZEROS_141  : slv141  := (others=>'0'); constant ZEROS_142  : slv142  := (others=>'0'); constant ZEROS_143  : slv143  := (others=>'0'); constant ZEROS_144  : slv144  := (others=>'0');
	constant ZEROS_145  : slv145  := (others=>'0'); constant ZEROS_146  : slv146  := (others=>'0'); constant ZEROS_147  : slv147  := (others=>'0'); constant ZEROS_148  : slv148  := (others=>'0');
	constant ZEROS_149  : slv149  := (others=>'0'); constant ZEROS_150  : slv150  := (others=>'0'); constant ZEROS_151  : slv151  := (others=>'0'); constant ZEROS_152  : slv152  := (others=>'0');
	constant ZEROS_153  : slv153  := (others=>'0'); constant ZEROS_154  : slv154  := (others=>'0'); constant ZEROS_155  : slv155  := (others=>'0'); constant ZEROS_156  : slv156  := (others=>'0');
	constant ZEROS_157  : slv157  := (others=>'0'); constant ZEROS_158  : slv158  := (others=>'0'); constant ZEROS_159  : slv159  := (others=>'0'); constant ZEROS_160  : slv160  := (others=>'0');
	constant ZEROS_161  : slv161  := (others=>'0'); constant ZEROS_162  : slv162  := (others=>'0'); constant ZEROS_163  : slv163  := (others=>'0'); constant ZEROS_164  : slv164  := (others=>'0');
	constant ZEROS_165  : slv165  := (others=>'0'); constant ZEROS_166  : slv166  := (others=>'0'); constant ZEROS_167  : slv167  := (others=>'0'); constant ZEROS_168  : slv168  := (others=>'0');
	constant ZEROS_169  : slv169  := (others=>'0'); constant ZEROS_170  : slv170  := (others=>'0'); constant ZEROS_171  : slv171  := (others=>'0'); constant ZEROS_172  : slv172  := (others=>'0');
	constant ZEROS_173  : slv173  := (others=>'0'); constant ZEROS_174  : slv174  := (others=>'0'); constant ZEROS_175  : slv175  := (others=>'0'); constant ZEROS_176  : slv176  := (others=>'0');
	constant ZEROS_177  : slv177  := (others=>'0'); constant ZEROS_178  : slv178  := (others=>'0'); constant ZEROS_179  : slv179  := (others=>'0'); constant ZEROS_180  : slv180  := (others=>'0');
	constant ZEROS_181  : slv181  := (others=>'0'); constant ZEROS_182  : slv182  := (others=>'0'); constant ZEROS_183  : slv183  := (others=>'0'); constant ZEROS_184  : slv184  := (others=>'0');
	constant ZEROS_185  : slv185  := (others=>'0'); constant ZEROS_186  : slv186  := (others=>'0'); constant ZEROS_187  : slv187  := (others=>'0'); constant ZEROS_188  : slv188  := (others=>'0');
	constant ZEROS_189  : slv189  := (others=>'0'); constant ZEROS_190  : slv190  := (others=>'0'); constant ZEROS_191  : slv191  := (others=>'0'); constant ZEROS_192  : slv192  := (others=>'0');
	constant ZEROS_193  : slv193  := (others=>'0'); constant ZEROS_194  : slv194  := (others=>'0'); constant ZEROS_195  : slv195  := (others=>'0'); constant ZEROS_196  : slv196  := (others=>'0');
	constant ZEROS_197  : slv197  := (others=>'0'); constant ZEROS_198  : slv198  := (others=>'0'); constant ZEROS_199  : slv199  := (others=>'0'); constant ZEROS_200  : slv200  := (others=>'0');
	constant ZEROS_201  : slv201  := (others=>'0'); constant ZEROS_202  : slv202  := (others=>'0'); constant ZEROS_203  : slv203  := (others=>'0'); constant ZEROS_204  : slv204  := (others=>'0');
	constant ZEROS_205  : slv205  := (others=>'0'); constant ZEROS_206  : slv206  := (others=>'0'); constant ZEROS_207  : slv207  := (others=>'0'); constant ZEROS_208  : slv208  := (others=>'0');
	constant ZEROS_209  : slv209  := (others=>'0'); constant ZEROS_210  : slv210  := (others=>'0'); constant ZEROS_211  : slv211  := (others=>'0'); constant ZEROS_212  : slv212  := (others=>'0');
	constant ZEROS_213  : slv213  := (others=>'0'); constant ZEROS_214  : slv214  := (others=>'0'); constant ZEROS_215  : slv215  := (others=>'0'); constant ZEROS_216  : slv216  := (others=>'0');
	constant ZEROS_217  : slv217  := (others=>'0'); constant ZEROS_218  : slv218  := (others=>'0'); constant ZEROS_219  : slv219  := (others=>'0'); constant ZEROS_220  : slv220  := (others=>'0');
	constant ZEROS_221  : slv221  := (others=>'0'); constant ZEROS_222  : slv222  := (others=>'0'); constant ZEROS_223  : slv223  := (others=>'0'); constant ZEROS_224  : slv224  := (others=>'0');
	constant ZEROS_225  : slv225  := (others=>'0'); constant ZEROS_226  : slv226  := (others=>'0'); constant ZEROS_227  : slv227  := (others=>'0'); constant ZEROS_228  : slv228  := (others=>'0');
	constant ZEROS_229  : slv229  := (others=>'0'); constant ZEROS_230  : slv230  := (others=>'0'); constant ZEROS_231  : slv231  := (others=>'0'); constant ZEROS_232  : slv232  := (others=>'0');
	constant ZEROS_233  : slv233  := (others=>'0'); constant ZEROS_234  : slv234  := (others=>'0'); constant ZEROS_235  : slv235  := (others=>'0'); constant ZEROS_236  : slv236  := (others=>'0');
	constant ZEROS_237  : slv237  := (others=>'0'); constant ZEROS_238  : slv238  := (others=>'0'); constant ZEROS_239  : slv239  := (others=>'0'); constant ZEROS_240  : slv240  := (others=>'0');
	constant ZEROS_241  : slv241  := (others=>'0'); constant ZEROS_242  : slv242  := (others=>'0'); constant ZEROS_243  : slv243  := (others=>'0'); constant ZEROS_244  : slv244  := (others=>'0');
	constant ZEROS_245  : slv245  := (others=>'0'); constant ZEROS_246  : slv246  := (others=>'0'); constant ZEROS_247  : slv247  := (others=>'0'); constant ZEROS_248  : slv248  := (others=>'0');
	constant ZEROS_249  : slv249  := (others=>'0'); constant ZEROS_250  : slv250  := (others=>'0'); constant ZEROS_251  : slv251  := (others=>'0'); constant ZEROS_252  : slv252  := (others=>'0');
	constant ZEROS_253  : slv253  := (others=>'0'); constant ZEROS_254  : slv254  := (others=>'0'); constant ZEROS_255  : slv255  := (others=>'0'); constant ZEROS_256  : slv256  := (others=>'0');
	constant ZEROS_257  : slv257  := (others=>'0'); constant ZEROS_258  : slv258  := (others=>'0'); constant ZEROS_259  : slv259  := (others=>'0'); constant ZEROS_260  : slv260  := (others=>'0');
	constant ZEROS_261  : slv261  := (others=>'0'); constant ZEROS_262  : slv262  := (others=>'0'); constant ZEROS_263  : slv263  := (others=>'0'); constant ZEROS_264  : slv264  := (others=>'0');
	constant ZEROS_265  : slv265  := (others=>'0'); constant ZEROS_266  : slv266  := (others=>'0'); constant ZEROS_267  : slv267  := (others=>'0'); constant ZEROS_268  : slv268  := (others=>'0');
	constant ZEROS_269  : slv269  := (others=>'0'); constant ZEROS_270  : slv270  := (others=>'0'); constant ZEROS_271  : slv271  := (others=>'0'); constant ZEROS_272  : slv272  := (others=>'0');
	constant ZEROS_273  : slv273  := (others=>'0'); constant ZEROS_274  : slv274  := (others=>'0'); constant ZEROS_275  : slv275  := (others=>'0'); constant ZEROS_276  : slv276  := (others=>'0');
	constant ZEROS_277  : slv277  := (others=>'0'); constant ZEROS_278  : slv278  := (others=>'0'); constant ZEROS_279  : slv279  := (others=>'0'); constant ZEROS_280  : slv280  := (others=>'0');
	constant ZEROS_281  : slv281  := (others=>'0'); constant ZEROS_282  : slv282  := (others=>'0'); constant ZEROS_283  : slv283  := (others=>'0'); constant ZEROS_284  : slv284  := (others=>'0');
	constant ZEROS_285  : slv285  := (others=>'0'); constant ZEROS_286  : slv286  := (others=>'0'); constant ZEROS_287  : slv287  := (others=>'0'); constant ZEROS_288  : slv288  := (others=>'0');
	constant ZEROS_289  : slv289  := (others=>'0'); constant ZEROS_290  : slv290  := (others=>'0'); constant ZEROS_291  : slv291  := (others=>'0'); constant ZEROS_292  : slv292  := (others=>'0');
	constant ZEROS_293  : slv293  := (others=>'0'); constant ZEROS_294  : slv294  := (others=>'0'); constant ZEROS_295  : slv295  := (others=>'0'); constant ZEROS_296  : slv296  := (others=>'0');
	constant ZEROS_297  : slv297  := (others=>'0'); constant ZEROS_298  : slv298  := (others=>'0'); constant ZEROS_299  : slv299  := (others=>'0'); constant ZEROS_300  : slv300  := (others=>'0');
	constant ZEROS_301  : slv301  := (others=>'0'); constant ZEROS_302  : slv302  := (others=>'0'); constant ZEROS_303  : slv303  := (others=>'0'); constant ZEROS_304  : slv304  := (others=>'0');
	constant ZEROS_305  : slv305  := (others=>'0'); constant ZEROS_306  : slv306  := (others=>'0'); constant ZEROS_307  : slv307  := (others=>'0'); constant ZEROS_308  : slv308  := (others=>'0');
	constant ZEROS_309  : slv309  := (others=>'0'); constant ZEROS_310  : slv310  := (others=>'0'); constant ZEROS_311  : slv311  := (others=>'0'); constant ZEROS_312  : slv312  := (others=>'0');
	constant ZEROS_313  : slv313  := (others=>'0'); constant ZEROS_314  : slv314  := (others=>'0'); constant ZEROS_315  : slv315  := (others=>'0'); constant ZEROS_316  : slv316  := (others=>'0');
	constant ZEROS_317  : slv317  := (others=>'0'); constant ZEROS_318  : slv318  := (others=>'0'); constant ZEROS_319  : slv319  := (others=>'0'); constant ZEROS_320  : slv320  := (others=>'0');
	constant ZEROS_321  : slv321  := (others=>'0'); constant ZEROS_322  : slv322  := (others=>'0'); constant ZEROS_323  : slv323  := (others=>'0'); constant ZEROS_324  : slv324  := (others=>'0');
	constant ZEROS_325  : slv325  := (others=>'0'); constant ZEROS_326  : slv326  := (others=>'0'); constant ZEROS_327  : slv327  := (others=>'0'); constant ZEROS_328  : slv328  := (others=>'0');
	constant ZEROS_329  : slv329  := (others=>'0'); constant ZEROS_330  : slv330  := (others=>'0'); constant ZEROS_331  : slv331  := (others=>'0'); constant ZEROS_332  : slv332  := (others=>'0');
	constant ZEROS_333  : slv333  := (others=>'0'); constant ZEROS_334  : slv334  := (others=>'0'); constant ZEROS_335  : slv335  := (others=>'0'); constant ZEROS_336  : slv336  := (others=>'0');
	constant ZEROS_337  : slv337  := (others=>'0'); constant ZEROS_338  : slv338  := (others=>'0'); constant ZEROS_339  : slv339  := (others=>'0'); constant ZEROS_340  : slv340  := (others=>'0');
	constant ZEROS_341  : slv341  := (others=>'0'); constant ZEROS_342  : slv342  := (others=>'0'); constant ZEROS_343  : slv343  := (others=>'0'); constant ZEROS_344  : slv344  := (others=>'0');
	constant ZEROS_345  : slv345  := (others=>'0'); constant ZEROS_346  : slv346  := (others=>'0'); constant ZEROS_347  : slv347  := (others=>'0'); constant ZEROS_348  : slv348  := (others=>'0');
	constant ZEROS_349  : slv349  := (others=>'0'); constant ZEROS_350  : slv350  := (others=>'0'); constant ZEROS_351  : slv351  := (others=>'0'); constant ZEROS_352  : slv352  := (others=>'0');
	constant ZEROS_353  : slv353  := (others=>'0'); constant ZEROS_354  : slv354  := (others=>'0'); constant ZEROS_355  : slv355  := (others=>'0'); constant ZEROS_356  : slv356  := (others=>'0');
	constant ZEROS_357  : slv357  := (others=>'0'); constant ZEROS_358  : slv358  := (others=>'0'); constant ZEROS_359  : slv359  := (others=>'0'); constant ZEROS_360  : slv360  := (others=>'0');
	constant ZEROS_361  : slv361  := (others=>'0'); constant ZEROS_362  : slv362  := (others=>'0'); constant ZEROS_363  : slv363  := (others=>'0'); constant ZEROS_364  : slv364  := (others=>'0');
	constant ZEROS_365  : slv365  := (others=>'0'); constant ZEROS_366  : slv366  := (others=>'0'); constant ZEROS_367  : slv367  := (others=>'0'); constant ZEROS_368  : slv368  := (others=>'0');
	constant ZEROS_369  : slv369  := (others=>'0'); constant ZEROS_370  : slv370  := (others=>'0'); constant ZEROS_371  : slv371  := (others=>'0'); constant ZEROS_372  : slv372  := (others=>'0');
	constant ZEROS_373  : slv373  := (others=>'0'); constant ZEROS_374  : slv374  := (others=>'0'); constant ZEROS_375  : slv375  := (others=>'0'); constant ZEROS_376  : slv376  := (others=>'0');
	constant ZEROS_377  : slv377  := (others=>'0'); constant ZEROS_378  : slv378  := (others=>'0'); constant ZEROS_379  : slv379  := (others=>'0'); constant ZEROS_380  : slv380  := (others=>'0');
	constant ZEROS_381  : slv381  := (others=>'0'); constant ZEROS_382  : slv382  := (others=>'0'); constant ZEROS_383  : slv383  := (others=>'0'); constant ZEROS_384  : slv384  := (others=>'0');
	constant ZEROS_385  : slv385  := (others=>'0'); constant ZEROS_386  : slv386  := (others=>'0'); constant ZEROS_387  : slv387  := (others=>'0'); constant ZEROS_388  : slv388  := (others=>'0');
	constant ZEROS_389  : slv389  := (others=>'0'); constant ZEROS_390  : slv390  := (others=>'0'); constant ZEROS_391  : slv391  := (others=>'0'); constant ZEROS_392  : slv392  := (others=>'0');
	constant ZEROS_393  : slv393  := (others=>'0'); constant ZEROS_394  : slv394  := (others=>'0'); constant ZEROS_395  : slv395  := (others=>'0'); constant ZEROS_396  : slv396  := (others=>'0');
	constant ZEROS_397  : slv397  := (others=>'0'); constant ZEROS_398  : slv398  := (others=>'0'); constant ZEROS_399  : slv399  := (others=>'0'); constant ZEROS_400  : slv400  := (others=>'0');
	constant ZEROS_401  : slv401  := (others=>'0'); constant ZEROS_402  : slv402  := (others=>'0'); constant ZEROS_403  : slv403  := (others=>'0'); constant ZEROS_404  : slv404  := (others=>'0');
	constant ZEROS_405  : slv405  := (others=>'0'); constant ZEROS_406  : slv406  := (others=>'0'); constant ZEROS_407  : slv407  := (others=>'0'); constant ZEROS_408  : slv408  := (others=>'0');
	constant ZEROS_409  : slv409  := (others=>'0'); constant ZEROS_410  : slv410  := (others=>'0'); constant ZEROS_411  : slv411  := (others=>'0'); constant ZEROS_412  : slv412  := (others=>'0');
	constant ZEROS_413  : slv413  := (others=>'0'); constant ZEROS_414  : slv414  := (others=>'0'); constant ZEROS_415  : slv415  := (others=>'0'); constant ZEROS_416  : slv416  := (others=>'0');
	constant ZEROS_417  : slv417  := (others=>'0'); constant ZEROS_418  : slv418  := (others=>'0'); constant ZEROS_419  : slv419  := (others=>'0'); constant ZEROS_420  : slv420  := (others=>'0');
	constant ZEROS_421  : slv421  := (others=>'0'); constant ZEROS_422  : slv422  := (others=>'0'); constant ZEROS_423  : slv423  := (others=>'0'); constant ZEROS_424  : slv424  := (others=>'0');
	constant ZEROS_425  : slv425  := (others=>'0'); constant ZEROS_426  : slv426  := (others=>'0'); constant ZEROS_427  : slv427  := (others=>'0'); constant ZEROS_428  : slv428  := (others=>'0');
	constant ZEROS_429  : slv429  := (others=>'0'); constant ZEROS_430  : slv430  := (others=>'0'); constant ZEROS_431  : slv431  := (others=>'0'); constant ZEROS_432  : slv432  := (others=>'0');
	constant ZEROS_433  : slv433  := (others=>'0'); constant ZEROS_434  : slv434  := (others=>'0'); constant ZEROS_435  : slv435  := (others=>'0'); constant ZEROS_436  : slv436  := (others=>'0');
	constant ZEROS_437  : slv437  := (others=>'0'); constant ZEROS_438  : slv438  := (others=>'0'); constant ZEROS_439  : slv439  := (others=>'0'); constant ZEROS_440  : slv440  := (others=>'0');
	constant ZEROS_441  : slv441  := (others=>'0'); constant ZEROS_442  : slv442  := (others=>'0'); constant ZEROS_443  : slv443  := (others=>'0'); constant ZEROS_444  : slv444  := (others=>'0');
	constant ZEROS_445  : slv445  := (others=>'0'); constant ZEROS_446  : slv446  := (others=>'0'); constant ZEROS_447  : slv447  := (others=>'0'); constant ZEROS_448  : slv448  := (others=>'0');
	constant ZEROS_449  : slv449  := (others=>'0'); constant ZEROS_450  : slv450  := (others=>'0'); constant ZEROS_451  : slv451  := (others=>'0'); constant ZEROS_452  : slv452  := (others=>'0');
	constant ZEROS_453  : slv453  := (others=>'0'); constant ZEROS_454  : slv454  := (others=>'0'); constant ZEROS_455  : slv455  := (others=>'0'); constant ZEROS_456  : slv456  := (others=>'0');
	constant ZEROS_457  : slv457  := (others=>'0'); constant ZEROS_458  : slv458  := (others=>'0'); constant ZEROS_459  : slv459  := (others=>'0'); constant ZEROS_460  : slv460  := (others=>'0');
	constant ZEROS_461  : slv461  := (others=>'0'); constant ZEROS_462  : slv462  := (others=>'0'); constant ZEROS_463  : slv463  := (others=>'0'); constant ZEROS_464  : slv464  := (others=>'0');
	constant ZEROS_465  : slv465  := (others=>'0'); constant ZEROS_466  : slv466  := (others=>'0'); constant ZEROS_467  : slv467  := (others=>'0'); constant ZEROS_468  : slv468  := (others=>'0');
	constant ZEROS_469  : slv469  := (others=>'0'); constant ZEROS_470  : slv470  := (others=>'0'); constant ZEROS_471  : slv471  := (others=>'0'); constant ZEROS_472  : slv472  := (others=>'0');
	constant ZEROS_473  : slv473  := (others=>'0'); constant ZEROS_474  : slv474  := (others=>'0'); constant ZEROS_475  : slv475  := (others=>'0'); constant ZEROS_476  : slv476  := (others=>'0');
	constant ZEROS_477  : slv477  := (others=>'0'); constant ZEROS_478  : slv478  := (others=>'0'); constant ZEROS_479  : slv479  := (others=>'0'); constant ZEROS_480  : slv480  := (others=>'0');
	constant ZEROS_481  : slv481  := (others=>'0'); constant ZEROS_482  : slv482  := (others=>'0'); constant ZEROS_483  : slv483  := (others=>'0'); constant ZEROS_484  : slv484  := (others=>'0');
	constant ZEROS_485  : slv485  := (others=>'0'); constant ZEROS_486  : slv486  := (others=>'0'); constant ZEROS_487  : slv487  := (others=>'0'); constant ZEROS_488  : slv488  := (others=>'0');
	constant ZEROS_489  : slv489  := (others=>'0'); constant ZEROS_490  : slv490  := (others=>'0'); constant ZEROS_491  : slv491  := (others=>'0'); constant ZEROS_492  : slv492  := (others=>'0');
	constant ZEROS_493  : slv493  := (others=>'0'); constant ZEROS_494  : slv494  := (others=>'0'); constant ZEROS_495  : slv495  := (others=>'0'); constant ZEROS_496  : slv496  := (others=>'0');
	constant ZEROS_497  : slv497  := (others=>'0'); constant ZEROS_498  : slv498  := (others=>'0'); constant ZEROS_499  : slv499  := (others=>'0'); constant ZEROS_500  : slv500  := (others=>'0');
	constant ZEROS_501  : slv501  := (others=>'0'); constant ZEROS_502  : slv502  := (others=>'0'); constant ZEROS_503  : slv503  := (others=>'0'); constant ZEROS_504  : slv504  := (others=>'0');
	constant ZEROS_505  : slv505  := (others=>'0'); constant ZEROS_506  : slv506  := (others=>'0'); constant ZEROS_507  : slv507  := (others=>'0'); constant ZEROS_508  : slv508  := (others=>'0');
	constant ZEROS_509  : slv509  := (others=>'0'); constant ZEROS_510  : slv510  := (others=>'0'); constant ZEROS_511  : slv511  := (others=>'0'); constant ZEROS_512  : slv512  := (others=>'0');
	constant ZEROS_513  : slv513  := (others=>'0'); constant ZEROS_514  : slv514  := (others=>'0'); constant ZEROS_515  : slv515  := (others=>'0'); constant ZEROS_516  : slv516  := (others=>'0');
	constant ZEROS_517  : slv517  := (others=>'0'); constant ZEROS_518  : slv518  := (others=>'0'); constant ZEROS_519  : slv519  := (others=>'0'); constant ZEROS_520  : slv520  := (others=>'0');
	constant ZEROS_521  : slv521  := (others=>'0'); constant ZEROS_522  : slv522  := (others=>'0'); constant ZEROS_523  : slv523  := (others=>'0'); constant ZEROS_524  : slv524  := (others=>'0');
	constant ZEROS_525  : slv525  := (others=>'0'); constant ZEROS_526  : slv526  := (others=>'0'); constant ZEROS_527  : slv527  := (others=>'0'); constant ZEROS_528  : slv528  := (others=>'0');
	constant ZEROS_529  : slv529  := (others=>'0'); constant ZEROS_530  : slv530  := (others=>'0'); constant ZEROS_531  : slv531  := (others=>'0'); constant ZEROS_532  : slv532  := (others=>'0');
	constant ZEROS_533  : slv533  := (others=>'0'); constant ZEROS_534  : slv534  := (others=>'0'); constant ZEROS_535  : slv535  := (others=>'0'); constant ZEROS_536  : slv536  := (others=>'0');
	constant ZEROS_537  : slv537  := (others=>'0'); constant ZEROS_538  : slv538  := (others=>'0'); constant ZEROS_539  : slv539  := (others=>'0'); constant ZEROS_540  : slv540  := (others=>'0');
	constant ZEROS_541  : slv541  := (others=>'0'); constant ZEROS_542  : slv542  := (others=>'0'); constant ZEROS_543  : slv543  := (others=>'0'); constant ZEROS_544  : slv544  := (others=>'0');
	constant ZEROS_545  : slv545  := (others=>'0'); constant ZEROS_546  : slv546  := (others=>'0'); constant ZEROS_547  : slv547  := (others=>'0'); constant ZEROS_548  : slv548  := (others=>'0');
	constant ZEROS_549  : slv549  := (others=>'0'); constant ZEROS_550  : slv550  := (others=>'0'); constant ZEROS_551  : slv551  := (others=>'0'); constant ZEROS_552  : slv552  := (others=>'0');
	constant ZEROS_553  : slv553  := (others=>'0'); constant ZEROS_554  : slv554  := (others=>'0'); constant ZEROS_555  : slv555  := (others=>'0'); constant ZEROS_556  : slv556  := (others=>'0');
	constant ZEROS_557  : slv557  := (others=>'0'); constant ZEROS_558  : slv558  := (others=>'0'); constant ZEROS_559  : slv559  := (others=>'0'); constant ZEROS_560  : slv560  := (others=>'0');
	constant ZEROS_561  : slv561  := (others=>'0'); constant ZEROS_562  : slv562  := (others=>'0'); constant ZEROS_563  : slv563  := (others=>'0'); constant ZEROS_564  : slv564  := (others=>'0');
	constant ZEROS_565  : slv565  := (others=>'0'); constant ZEROS_566  : slv566  := (others=>'0'); constant ZEROS_567  : slv567  := (others=>'0'); constant ZEROS_568  : slv568  := (others=>'0');
	constant ZEROS_569  : slv569  := (others=>'0'); constant ZEROS_570  : slv570  := (others=>'0'); constant ZEROS_571  : slv571  := (others=>'0'); constant ZEROS_572  : slv572  := (others=>'0');
	constant ZEROS_573  : slv573  := (others=>'0'); constant ZEROS_574  : slv574  := (others=>'0'); constant ZEROS_575  : slv575  := (others=>'0'); constant ZEROS_576  : slv576  := (others=>'0');
	constant ZEROS_577  : slv577  := (others=>'0'); constant ZEROS_578  : slv578  := (others=>'0'); constant ZEROS_579  : slv579  := (others=>'0'); constant ZEROS_580  : slv580  := (others=>'0');
	constant ZEROS_581  : slv581  := (others=>'0'); constant ZEROS_582  : slv582  := (others=>'0'); constant ZEROS_583  : slv583  := (others=>'0'); constant ZEROS_584  : slv584  := (others=>'0');
	constant ZEROS_585  : slv585  := (others=>'0'); constant ZEROS_586  : slv586  := (others=>'0'); constant ZEROS_587  : slv587  := (others=>'0'); constant ZEROS_588  : slv588  := (others=>'0');
	constant ZEROS_589  : slv589  := (others=>'0'); constant ZEROS_590  : slv590  := (others=>'0'); constant ZEROS_591  : slv591  := (others=>'0'); constant ZEROS_592  : slv592  := (others=>'0');
	constant ZEROS_593  : slv593  := (others=>'0'); constant ZEROS_594  : slv594  := (others=>'0'); constant ZEROS_595  : slv595  := (others=>'0'); constant ZEROS_596  : slv596  := (others=>'0');
	constant ZEROS_597  : slv597  := (others=>'0'); constant ZEROS_598  : slv598  := (others=>'0'); constant ZEROS_599  : slv599  := (others=>'0'); constant ZEROS_600  : slv600  := (others=>'0');
	constant ZEROS_601  : slv601  := (others=>'0'); constant ZEROS_602  : slv602  := (others=>'0'); constant ZEROS_603  : slv603  := (others=>'0'); constant ZEROS_604  : slv604  := (others=>'0');
	constant ZEROS_605  : slv605  := (others=>'0'); constant ZEROS_606  : slv606  := (others=>'0'); constant ZEROS_607  : slv607  := (others=>'0'); constant ZEROS_608  : slv608  := (others=>'0');
	constant ZEROS_609  : slv609  := (others=>'0'); constant ZEROS_610  : slv610  := (others=>'0'); constant ZEROS_611  : slv611  := (others=>'0'); constant ZEROS_612  : slv612  := (others=>'0');
	constant ZEROS_613  : slv613  := (others=>'0'); constant ZEROS_614  : slv614  := (others=>'0'); constant ZEROS_615  : slv615  := (others=>'0'); constant ZEROS_616  : slv616  := (others=>'0');
	constant ZEROS_617  : slv617  := (others=>'0'); constant ZEROS_618  : slv618  := (others=>'0'); constant ZEROS_619  : slv619  := (others=>'0'); constant ZEROS_620  : slv620  := (others=>'0');
	constant ZEROS_621  : slv621  := (others=>'0'); constant ZEROS_622  : slv622  := (others=>'0'); constant ZEROS_623  : slv623  := (others=>'0'); constant ZEROS_624  : slv624  := (others=>'0');
	constant ZEROS_625  : slv625  := (others=>'0'); constant ZEROS_626  : slv626  := (others=>'0'); constant ZEROS_627  : slv627  := (others=>'0'); constant ZEROS_628  : slv628  := (others=>'0');
	constant ZEROS_629  : slv629  := (others=>'0'); constant ZEROS_630  : slv630  := (others=>'0'); constant ZEROS_631  : slv631  := (others=>'0'); constant ZEROS_632  : slv632  := (others=>'0');
	constant ZEROS_633  : slv633  := (others=>'0'); constant ZEROS_634  : slv634  := (others=>'0'); constant ZEROS_635  : slv635  := (others=>'0'); constant ZEROS_636  : slv636  := (others=>'0');
	constant ZEROS_637  : slv637  := (others=>'0'); constant ZEROS_638  : slv638  := (others=>'0'); constant ZEROS_639  : slv639  := (others=>'0'); constant ZEROS_640  : slv640  := (others=>'0');
	constant ZEROS_641  : slv641  := (others=>'0'); constant ZEROS_642  : slv642  := (others=>'0'); constant ZEROS_643  : slv643  := (others=>'0'); constant ZEROS_644  : slv644  := (others=>'0');
	constant ZEROS_645  : slv645  := (others=>'0'); constant ZEROS_646  : slv646  := (others=>'0'); constant ZEROS_647  : slv647  := (others=>'0'); constant ZEROS_648  : slv648  := (others=>'0');
	constant ZEROS_649  : slv649  := (others=>'0'); constant ZEROS_650  : slv650  := (others=>'0'); constant ZEROS_651  : slv651  := (others=>'0'); constant ZEROS_652  : slv652  := (others=>'0');
	constant ZEROS_653  : slv653  := (others=>'0'); constant ZEROS_654  : slv654  := (others=>'0'); constant ZEROS_655  : slv655  := (others=>'0'); constant ZEROS_656  : slv656  := (others=>'0');
	constant ZEROS_657  : slv657  := (others=>'0'); constant ZEROS_658  : slv658  := (others=>'0'); constant ZEROS_659  : slv659  := (others=>'0'); constant ZEROS_660  : slv660  := (others=>'0');
	constant ZEROS_661  : slv661  := (others=>'0'); constant ZEROS_662  : slv662  := (others=>'0'); constant ZEROS_663  : slv663  := (others=>'0'); constant ZEROS_664  : slv664  := (others=>'0');
	constant ZEROS_665  : slv665  := (others=>'0'); constant ZEROS_666  : slv666  := (others=>'0'); constant ZEROS_667  : slv667  := (others=>'0'); constant ZEROS_668  : slv668  := (others=>'0');
	constant ZEROS_669  : slv669  := (others=>'0'); constant ZEROS_670  : slv670  := (others=>'0'); constant ZEROS_671  : slv671  := (others=>'0'); constant ZEROS_672  : slv672  := (others=>'0');
	constant ZEROS_673  : slv673  := (others=>'0'); constant ZEROS_674  : slv674  := (others=>'0'); constant ZEROS_675  : slv675  := (others=>'0'); constant ZEROS_676  : slv676  := (others=>'0');
	constant ZEROS_677  : slv677  := (others=>'0'); constant ZEROS_678  : slv678  := (others=>'0'); constant ZEROS_679  : slv679  := (others=>'0'); constant ZEROS_680  : slv680  := (others=>'0');
	constant ZEROS_681  : slv681  := (others=>'0'); constant ZEROS_682  : slv682  := (others=>'0'); constant ZEROS_683  : slv683  := (others=>'0'); constant ZEROS_684  : slv684  := (others=>'0');
	constant ZEROS_685  : slv685  := (others=>'0'); constant ZEROS_686  : slv686  := (others=>'0'); constant ZEROS_687  : slv687  := (others=>'0'); constant ZEROS_688  : slv688  := (others=>'0');
	constant ZEROS_689  : slv689  := (others=>'0'); constant ZEROS_690  : slv690  := (others=>'0'); constant ZEROS_691  : slv691  := (others=>'0'); constant ZEROS_692  : slv692  := (others=>'0');
	constant ZEROS_693  : slv693  := (others=>'0'); constant ZEROS_694  : slv694  := (others=>'0'); constant ZEROS_695  : slv695  := (others=>'0'); constant ZEROS_696  : slv696  := (others=>'0');
	constant ZEROS_697  : slv697  := (others=>'0'); constant ZEROS_698  : slv698  := (others=>'0'); constant ZEROS_699  : slv699  := (others=>'0'); constant ZEROS_700  : slv700  := (others=>'0');
	constant ZEROS_701  : slv701  := (others=>'0'); constant ZEROS_702  : slv702  := (others=>'0'); constant ZEROS_703  : slv703  := (others=>'0'); constant ZEROS_704  : slv704  := (others=>'0');
	constant ZEROS_705  : slv705  := (others=>'0'); constant ZEROS_706  : slv706  := (others=>'0'); constant ZEROS_707  : slv707  := (others=>'0'); constant ZEROS_708  : slv708  := (others=>'0');
	constant ZEROS_709  : slv709  := (others=>'0'); constant ZEROS_710  : slv710  := (others=>'0'); constant ZEROS_711  : slv711  := (others=>'0'); constant ZEROS_712  : slv712  := (others=>'0');
	constant ZEROS_713  : slv713  := (others=>'0'); constant ZEROS_714  : slv714  := (others=>'0'); constant ZEROS_715  : slv715  := (others=>'0'); constant ZEROS_716  : slv716  := (others=>'0');
	constant ZEROS_717  : slv717  := (others=>'0'); constant ZEROS_718  : slv718  := (others=>'0'); constant ZEROS_719  : slv719  := (others=>'0'); constant ZEROS_720  : slv720  := (others=>'0');
	constant ZEROS_721  : slv721  := (others=>'0'); constant ZEROS_722  : slv722  := (others=>'0'); constant ZEROS_723  : slv723  := (others=>'0'); constant ZEROS_724  : slv724  := (others=>'0');
	constant ZEROS_725  : slv725  := (others=>'0'); constant ZEROS_726  : slv726  := (others=>'0'); constant ZEROS_727  : slv727  := (others=>'0'); constant ZEROS_728  : slv728  := (others=>'0');
	constant ZEROS_729  : slv729  := (others=>'0'); constant ZEROS_730  : slv730  := (others=>'0'); constant ZEROS_731  : slv731  := (others=>'0'); constant ZEROS_732  : slv732  := (others=>'0');
	constant ZEROS_733  : slv733  := (others=>'0'); constant ZEROS_734  : slv734  := (others=>'0'); constant ZEROS_735  : slv735  := (others=>'0'); constant ZEROS_736  : slv736  := (others=>'0');
	constant ZEROS_737  : slv737  := (others=>'0'); constant ZEROS_738  : slv738  := (others=>'0'); constant ZEROS_739  : slv739  := (others=>'0'); constant ZEROS_740  : slv740  := (others=>'0');
	constant ZEROS_741  : slv741  := (others=>'0'); constant ZEROS_742  : slv742  := (others=>'0'); constant ZEROS_743  : slv743  := (others=>'0'); constant ZEROS_744  : slv744  := (others=>'0');
	constant ZEROS_745  : slv745  := (others=>'0'); constant ZEROS_746  : slv746  := (others=>'0'); constant ZEROS_747  : slv747  := (others=>'0'); constant ZEROS_748  : slv748  := (others=>'0');
	constant ZEROS_749  : slv749  := (others=>'0'); constant ZEROS_750  : slv750  := (others=>'0'); constant ZEROS_751  : slv751  := (others=>'0'); constant ZEROS_752  : slv752  := (others=>'0');
	constant ZEROS_753  : slv753  := (others=>'0'); constant ZEROS_754  : slv754  := (others=>'0'); constant ZEROS_755  : slv755  := (others=>'0'); constant ZEROS_756  : slv756  := (others=>'0');
	constant ZEROS_757  : slv757  := (others=>'0'); constant ZEROS_758  : slv758  := (others=>'0'); constant ZEROS_759  : slv759  := (others=>'0'); constant ZEROS_760  : slv760  := (others=>'0');
	constant ZEROS_761  : slv761  := (others=>'0'); constant ZEROS_762  : slv762  := (others=>'0'); constant ZEROS_763  : slv763  := (others=>'0'); constant ZEROS_764  : slv764  := (others=>'0');
	constant ZEROS_765  : slv765  := (others=>'0'); constant ZEROS_766  : slv766  := (others=>'0'); constant ZEROS_767  : slv767  := (others=>'0'); constant ZEROS_768  : slv768  := (others=>'0');
	constant ZEROS_769  : slv769  := (others=>'0'); constant ZEROS_770  : slv770  := (others=>'0'); constant ZEROS_771  : slv771  := (others=>'0'); constant ZEROS_772  : slv772  := (others=>'0');
	constant ZEROS_773  : slv773  := (others=>'0'); constant ZEROS_774  : slv774  := (others=>'0'); constant ZEROS_775  : slv775  := (others=>'0'); constant ZEROS_776  : slv776  := (others=>'0');
	constant ZEROS_777  : slv777  := (others=>'0'); constant ZEROS_778  : slv778  := (others=>'0'); constant ZEROS_779  : slv779  := (others=>'0'); constant ZEROS_780  : slv780  := (others=>'0');
	constant ZEROS_781  : slv781  := (others=>'0'); constant ZEROS_782  : slv782  := (others=>'0'); constant ZEROS_783  : slv783  := (others=>'0'); constant ZEROS_784  : slv784  := (others=>'0');
	constant ZEROS_785  : slv785  := (others=>'0'); constant ZEROS_786  : slv786  := (others=>'0'); constant ZEROS_787  : slv787  := (others=>'0'); constant ZEROS_788  : slv788  := (others=>'0');
	constant ZEROS_789  : slv789  := (others=>'0'); constant ZEROS_790  : slv790  := (others=>'0'); constant ZEROS_791  : slv791  := (others=>'0'); constant ZEROS_792  : slv792  := (others=>'0');
	constant ZEROS_793  : slv793  := (others=>'0'); constant ZEROS_794  : slv794  := (others=>'0'); constant ZEROS_795  : slv795  := (others=>'0'); constant ZEROS_796  : slv796  := (others=>'0');
	constant ZEROS_797  : slv797  := (others=>'0'); constant ZEROS_798  : slv798  := (others=>'0'); constant ZEROS_799  : slv799  := (others=>'0'); constant ZEROS_800  : slv800  := (others=>'0');
	constant ZEROS_801  : slv801  := (others=>'0'); constant ZEROS_802  : slv802  := (others=>'0'); constant ZEROS_803  : slv803  := (others=>'0'); constant ZEROS_804  : slv804  := (others=>'0');
	constant ZEROS_805  : slv805  := (others=>'0'); constant ZEROS_806  : slv806  := (others=>'0'); constant ZEROS_807  : slv807  := (others=>'0'); constant ZEROS_808  : slv808  := (others=>'0');
	constant ZEROS_809  : slv809  := (others=>'0'); constant ZEROS_810  : slv810  := (others=>'0'); constant ZEROS_811  : slv811  := (others=>'0'); constant ZEROS_812  : slv812  := (others=>'0');
	constant ZEROS_813  : slv813  := (others=>'0'); constant ZEROS_814  : slv814  := (others=>'0'); constant ZEROS_815  : slv815  := (others=>'0'); constant ZEROS_816  : slv816  := (others=>'0');
	constant ZEROS_817  : slv817  := (others=>'0'); constant ZEROS_818  : slv818  := (others=>'0'); constant ZEROS_819  : slv819  := (others=>'0'); constant ZEROS_820  : slv820  := (others=>'0');
	constant ZEROS_821  : slv821  := (others=>'0'); constant ZEROS_822  : slv822  := (others=>'0'); constant ZEROS_823  : slv823  := (others=>'0'); constant ZEROS_824  : slv824  := (others=>'0');
	constant ZEROS_825  : slv825  := (others=>'0'); constant ZEROS_826  : slv826  := (others=>'0'); constant ZEROS_827  : slv827  := (others=>'0'); constant ZEROS_828  : slv828  := (others=>'0');
	constant ZEROS_829  : slv829  := (others=>'0'); constant ZEROS_830  : slv830  := (others=>'0'); constant ZEROS_831  : slv831  := (others=>'0'); constant ZEROS_832  : slv832  := (others=>'0');
	constant ZEROS_833  : slv833  := (others=>'0'); constant ZEROS_834  : slv834  := (others=>'0'); constant ZEROS_835  : slv835  := (others=>'0'); constant ZEROS_836  : slv836  := (others=>'0');
	constant ZEROS_837  : slv837  := (others=>'0'); constant ZEROS_838  : slv838  := (others=>'0'); constant ZEROS_839  : slv839  := (others=>'0'); constant ZEROS_840  : slv840  := (others=>'0');
	constant ZEROS_841  : slv841  := (others=>'0'); constant ZEROS_842  : slv842  := (others=>'0'); constant ZEROS_843  : slv843  := (others=>'0'); constant ZEROS_844  : slv844  := (others=>'0');
	constant ZEROS_845  : slv845  := (others=>'0'); constant ZEROS_846  : slv846  := (others=>'0'); constant ZEROS_847  : slv847  := (others=>'0'); constant ZEROS_848  : slv848  := (others=>'0');
	constant ZEROS_849  : slv849  := (others=>'0'); constant ZEROS_850  : slv850  := (others=>'0'); constant ZEROS_851  : slv851  := (others=>'0'); constant ZEROS_852  : slv852  := (others=>'0');
	constant ZEROS_853  : slv853  := (others=>'0'); constant ZEROS_854  : slv854  := (others=>'0'); constant ZEROS_855  : slv855  := (others=>'0'); constant ZEROS_856  : slv856  := (others=>'0');
	constant ZEROS_857  : slv857  := (others=>'0'); constant ZEROS_858  : slv858  := (others=>'0'); constant ZEROS_859  : slv859  := (others=>'0'); constant ZEROS_860  : slv860  := (others=>'0');
	constant ZEROS_861  : slv861  := (others=>'0'); constant ZEROS_862  : slv862  := (others=>'0'); constant ZEROS_863  : slv863  := (others=>'0'); constant ZEROS_864  : slv864  := (others=>'0');
	constant ZEROS_865  : slv865  := (others=>'0'); constant ZEROS_866  : slv866  := (others=>'0'); constant ZEROS_867  : slv867  := (others=>'0'); constant ZEROS_868  : slv868  := (others=>'0');
	constant ZEROS_869  : slv869  := (others=>'0'); constant ZEROS_870  : slv870  := (others=>'0'); constant ZEROS_871  : slv871  := (others=>'0'); constant ZEROS_872  : slv872  := (others=>'0');
	constant ZEROS_873  : slv873  := (others=>'0'); constant ZEROS_874  : slv874  := (others=>'0'); constant ZEROS_875  : slv875  := (others=>'0'); constant ZEROS_876  : slv876  := (others=>'0');
	constant ZEROS_877  : slv877  := (others=>'0'); constant ZEROS_878  : slv878  := (others=>'0'); constant ZEROS_879  : slv879  := (others=>'0'); constant ZEROS_880  : slv880  := (others=>'0');
	constant ZEROS_881  : slv881  := (others=>'0'); constant ZEROS_882  : slv882  := (others=>'0'); constant ZEROS_883  : slv883  := (others=>'0'); constant ZEROS_884  : slv884  := (others=>'0');
	constant ZEROS_885  : slv885  := (others=>'0'); constant ZEROS_886  : slv886  := (others=>'0'); constant ZEROS_887  : slv887  := (others=>'0'); constant ZEROS_888  : slv888  := (others=>'0');
	constant ZEROS_889  : slv889  := (others=>'0'); constant ZEROS_890  : slv890  := (others=>'0'); constant ZEROS_891  : slv891  := (others=>'0'); constant ZEROS_892  : slv892  := (others=>'0');
	constant ZEROS_893  : slv893  := (others=>'0'); constant ZEROS_894  : slv894  := (others=>'0'); constant ZEROS_895  : slv895  := (others=>'0'); constant ZEROS_896  : slv896  := (others=>'0');
	constant ZEROS_897  : slv897  := (others=>'0'); constant ZEROS_898  : slv898  := (others=>'0'); constant ZEROS_899  : slv899  := (others=>'0'); constant ZEROS_900  : slv900  := (others=>'0');
	constant ZEROS_901  : slv901  := (others=>'0'); constant ZEROS_902  : slv902  := (others=>'0'); constant ZEROS_903  : slv903  := (others=>'0'); constant ZEROS_904  : slv904  := (others=>'0');
	constant ZEROS_905  : slv905  := (others=>'0'); constant ZEROS_906  : slv906  := (others=>'0'); constant ZEROS_907  : slv907  := (others=>'0'); constant ZEROS_908  : slv908  := (others=>'0');
	constant ZEROS_909  : slv909  := (others=>'0'); constant ZEROS_910  : slv910  := (others=>'0'); constant ZEROS_911  : slv911  := (others=>'0'); constant ZEROS_912  : slv912  := (others=>'0');
	constant ZEROS_913  : slv913  := (others=>'0'); constant ZEROS_914  : slv914  := (others=>'0'); constant ZEROS_915  : slv915  := (others=>'0'); constant ZEROS_916  : slv916  := (others=>'0');
	constant ZEROS_917  : slv917  := (others=>'0'); constant ZEROS_918  : slv918  := (others=>'0'); constant ZEROS_919  : slv919  := (others=>'0'); constant ZEROS_920  : slv920  := (others=>'0');
	constant ZEROS_921  : slv921  := (others=>'0'); constant ZEROS_922  : slv922  := (others=>'0'); constant ZEROS_923  : slv923  := (others=>'0'); constant ZEROS_924  : slv924  := (others=>'0');
	constant ZEROS_925  : slv925  := (others=>'0'); constant ZEROS_926  : slv926  := (others=>'0'); constant ZEROS_927  : slv927  := (others=>'0'); constant ZEROS_928  : slv928  := (others=>'0');
	constant ZEROS_929  : slv929  := (others=>'0'); constant ZEROS_930  : slv930  := (others=>'0'); constant ZEROS_931  : slv931  := (others=>'0'); constant ZEROS_932  : slv932  := (others=>'0');
	constant ZEROS_933  : slv933  := (others=>'0'); constant ZEROS_934  : slv934  := (others=>'0'); constant ZEROS_935  : slv935  := (others=>'0'); constant ZEROS_936  : slv936  := (others=>'0');
	constant ZEROS_937  : slv937  := (others=>'0'); constant ZEROS_938  : slv938  := (others=>'0'); constant ZEROS_939  : slv939  := (others=>'0'); constant ZEROS_940  : slv940  := (others=>'0');
	constant ZEROS_941  : slv941  := (others=>'0'); constant ZEROS_942  : slv942  := (others=>'0'); constant ZEROS_943  : slv943  := (others=>'0'); constant ZEROS_944  : slv944  := (others=>'0');
	constant ZEROS_945  : slv945  := (others=>'0'); constant ZEROS_946  : slv946  := (others=>'0'); constant ZEROS_947  : slv947  := (others=>'0'); constant ZEROS_948  : slv948  := (others=>'0');
	constant ZEROS_949  : slv949  := (others=>'0'); constant ZEROS_950  : slv950  := (others=>'0'); constant ZEROS_951  : slv951  := (others=>'0'); constant ZEROS_952  : slv952  := (others=>'0');
	constant ZEROS_953  : slv953  := (others=>'0'); constant ZEROS_954  : slv954  := (others=>'0'); constant ZEROS_955  : slv955  := (others=>'0'); constant ZEROS_956  : slv956  := (others=>'0');
	constant ZEROS_957  : slv957  := (others=>'0'); constant ZEROS_958  : slv958  := (others=>'0'); constant ZEROS_959  : slv959  := (others=>'0'); constant ZEROS_960  : slv960  := (others=>'0');
	constant ZEROS_961  : slv961  := (others=>'0'); constant ZEROS_962  : slv962  := (others=>'0'); constant ZEROS_963  : slv963  := (others=>'0'); constant ZEROS_964  : slv964  := (others=>'0');
	constant ZEROS_965  : slv965  := (others=>'0'); constant ZEROS_966  : slv966  := (others=>'0'); constant ZEROS_967  : slv967  := (others=>'0'); constant ZEROS_968  : slv968  := (others=>'0');
	constant ZEROS_969  : slv969  := (others=>'0'); constant ZEROS_970  : slv970  := (others=>'0'); constant ZEROS_971  : slv971  := (others=>'0'); constant ZEROS_972  : slv972  := (others=>'0');
	constant ZEROS_973  : slv973  := (others=>'0'); constant ZEROS_974  : slv974  := (others=>'0'); constant ZEROS_975  : slv975  := (others=>'0'); constant ZEROS_976  : slv976  := (others=>'0');
	constant ZEROS_977  : slv977  := (others=>'0'); constant ZEROS_978  : slv978  := (others=>'0'); constant ZEROS_979  : slv979  := (others=>'0'); constant ZEROS_980  : slv980  := (others=>'0');
	constant ZEROS_981  : slv981  := (others=>'0'); constant ZEROS_982  : slv982  := (others=>'0'); constant ZEROS_983  : slv983  := (others=>'0'); constant ZEROS_984  : slv984  := (others=>'0');
	constant ZEROS_985  : slv985  := (others=>'0'); constant ZEROS_986  : slv986  := (others=>'0'); constant ZEROS_987  : slv987  := (others=>'0'); constant ZEROS_988  : slv988  := (others=>'0');
	constant ZEROS_989  : slv989  := (others=>'0'); constant ZEROS_990  : slv990  := (others=>'0'); constant ZEROS_991  : slv991  := (others=>'0'); constant ZEROS_992  : slv992  := (others=>'0');
	constant ZEROS_993  : slv993  := (others=>'0'); constant ZEROS_994  : slv994  := (others=>'0'); constant ZEROS_995  : slv995  := (others=>'0'); constant ZEROS_996  : slv996  := (others=>'0');
	constant ZEROS_997  : slv997  := (others=>'0'); constant ZEROS_998  : slv998  := (others=>'0'); constant ZEROS_999  : slv999  := (others=>'0'); constant ZEROS_1000 : slv1000 := (others=>'0');
	constant ZEROS_1001 : slv1001 := (others=>'0'); constant ZEROS_1002 : slv1002 := (others=>'0'); constant ZEROS_1003 : slv1003 := (others=>'0'); constant ZEROS_1004 : slv1004 := (others=>'0');
	constant ZEROS_1005 : slv1005 := (others=>'0'); constant ZEROS_1006 : slv1006 := (others=>'0'); constant ZEROS_1007 : slv1007 := (others=>'0'); constant ZEROS_1008 : slv1008 := (others=>'0');
	constant ZEROS_1009 : slv1009 := (others=>'0'); constant ZEROS_1010 : slv1010 := (others=>'0'); constant ZEROS_1011 : slv1011 := (others=>'0'); constant ZEROS_1012 : slv1012 := (others=>'0');
	constant ZEROS_1013 : slv1013 := (others=>'0'); constant ZEROS_1014 : slv1014 := (others=>'0'); constant ZEROS_1015 : slv1015 := (others=>'0'); constant ZEROS_1016 : slv1016 := (others=>'0');
	constant ZEROS_1017 : slv1017 := (others=>'0'); constant ZEROS_1018 : slv1018 := (others=>'0'); constant ZEROS_1019 : slv1019 := (others=>'0'); constant ZEROS_1020 : slv1020 := (others=>'0');
	constant ZEROS_1021 : slv1021 := (others=>'0'); constant ZEROS_1022 : slv1022 := (others=>'0'); constant ZEROS_1023 : slv1023 := (others=>'0'); constant ZEROS_1024 : slv1024 := (others=>'0');
--**************************************************************************************************************************************************************
-- ONE
--**************************************************************************************************************************************************************
	constant ONES      : slv(1023 downto 0) := (others=>'1');
	constant ONES_1    : slv1    := (others=>'1'); constant ONES_2    : slv2    := (others=>'1'); constant ONES_3    : slv3    := (others=>'1'); constant ONES_4    : slv4    := (others=>'1');
	constant ONES_5    : slv5    := (others=>'1'); constant ONES_6    : slv6    := (others=>'1'); constant ONES_7    : slv7    := (others=>'1'); constant ONES_8    : slv8    := (others=>'1');
	constant ONES_9    : slv9    := (others=>'1'); constant ONES_10   : slv10   := (others=>'1'); constant ONES_11   : slv11   := (others=>'1'); constant ONES_12   : slv12   := (others=>'1');
	constant ONES_13   : slv13   := (others=>'1'); constant ONES_14   : slv14   := (others=>'1'); constant ONES_15   : slv15   := (others=>'1'); constant ONES_16   : slv16   := (others=>'1');
	constant ONES_17   : slv17   := (others=>'1'); constant ONES_18   : slv18   := (others=>'1'); constant ONES_19   : slv19   := (others=>'1'); constant ONES_20   : slv20   := (others=>'1');
	constant ONES_21   : slv21   := (others=>'1'); constant ONES_22   : slv22   := (others=>'1'); constant ONES_23   : slv23   := (others=>'1'); constant ONES_24   : slv24   := (others=>'1');
	constant ONES_25   : slv25   := (others=>'1'); constant ONES_26   : slv26   := (others=>'1'); constant ONES_27   : slv27   := (others=>'1'); constant ONES_28   : slv28   := (others=>'1');
	constant ONES_29   : slv29   := (others=>'1'); constant ONES_30   : slv30   := (others=>'1'); constant ONES_31   : slv31   := (others=>'1'); constant ONES_32   : slv32   := (others=>'1');
	constant ONES_33   : slv33   := (others=>'1'); constant ONES_34   : slv34   := (others=>'1'); constant ONES_35   : slv35   := (others=>'1'); constant ONES_36   : slv36   := (others=>'1');
	constant ONES_37   : slv37   := (others=>'1'); constant ONES_38   : slv38   := (others=>'1'); constant ONES_39   : slv39   := (others=>'1'); constant ONES_40   : slv40   := (others=>'1');
	constant ONES_41   : slv41   := (others=>'1'); constant ONES_42   : slv42   := (others=>'1'); constant ONES_43   : slv43   := (others=>'1'); constant ONES_44   : slv44   := (others=>'1');
	constant ONES_45   : slv45   := (others=>'1'); constant ONES_46   : slv46   := (others=>'1'); constant ONES_47   : slv47   := (others=>'1'); constant ONES_48   : slv48   := (others=>'1');
	constant ONES_49   : slv49   := (others=>'1'); constant ONES_50   : slv50   := (others=>'1'); constant ONES_51   : slv51   := (others=>'1'); constant ONES_52   : slv52   := (others=>'1');
	constant ONES_53   : slv53   := (others=>'1'); constant ONES_54   : slv54   := (others=>'1'); constant ONES_55   : slv55   := (others=>'1'); constant ONES_56   : slv56   := (others=>'1');
	constant ONES_57   : slv57   := (others=>'1'); constant ONES_58   : slv58   := (others=>'1'); constant ONES_59   : slv59   := (others=>'1'); constant ONES_60   : slv60   := (others=>'1');
	constant ONES_61   : slv61   := (others=>'1'); constant ONES_62   : slv62   := (others=>'1'); constant ONES_63   : slv63   := (others=>'1'); constant ONES_64   : slv64   := (others=>'1');
	constant ONES_65   : slv65   := (others=>'1'); constant ONES_66   : slv66   := (others=>'1'); constant ONES_67   : slv67   := (others=>'1'); constant ONES_68   : slv68   := (others=>'1');
	constant ONES_69   : slv69   := (others=>'1'); constant ONES_70   : slv70   := (others=>'1'); constant ONES_71   : slv71   := (others=>'1'); constant ONES_72   : slv72   := (others=>'1');
	constant ONES_73   : slv73   := (others=>'1'); constant ONES_74   : slv74   := (others=>'1'); constant ONES_75   : slv75   := (others=>'1'); constant ONES_76   : slv76   := (others=>'1');
	constant ONES_77   : slv77   := (others=>'1'); constant ONES_78   : slv78   := (others=>'1'); constant ONES_79   : slv79   := (others=>'1'); constant ONES_80   : slv80   := (others=>'1');
	constant ONES_81   : slv81   := (others=>'1'); constant ONES_82   : slv82   := (others=>'1'); constant ONES_83   : slv83   := (others=>'1'); constant ONES_84   : slv84   := (others=>'1');
	constant ONES_85   : slv85   := (others=>'1'); constant ONES_86   : slv86   := (others=>'1'); constant ONES_87   : slv87   := (others=>'1'); constant ONES_88   : slv88   := (others=>'1');
	constant ONES_89   : slv89   := (others=>'1'); constant ONES_90   : slv90   := (others=>'1'); constant ONES_91   : slv91   := (others=>'1'); constant ONES_92   : slv92   := (others=>'1');
	constant ONES_93   : slv93   := (others=>'1'); constant ONES_94   : slv94   := (others=>'1'); constant ONES_95   : slv95   := (others=>'1'); constant ONES_96   : slv96   := (others=>'1');
	constant ONES_97   : slv97   := (others=>'1'); constant ONES_98   : slv98   := (others=>'1'); constant ONES_99   : slv99   := (others=>'1'); constant ONES_100  : slv100  := (others=>'1');
	constant ONES_101  : slv101  := (others=>'1'); constant ONES_102  : slv102  := (others=>'1'); constant ONES_103  : slv103  := (others=>'1'); constant ONES_104  : slv104  := (others=>'1');
	constant ONES_105  : slv105  := (others=>'1'); constant ONES_106  : slv106  := (others=>'1'); constant ONES_107  : slv107  := (others=>'1'); constant ONES_108  : slv108  := (others=>'1');
	constant ONES_109  : slv109  := (others=>'1'); constant ONES_110  : slv110  := (others=>'1'); constant ONES_111  : slv111  := (others=>'1'); constant ONES_112  : slv112  := (others=>'1');
	constant ONES_113  : slv113  := (others=>'1'); constant ONES_114  : slv114  := (others=>'1'); constant ONES_115  : slv115  := (others=>'1'); constant ONES_116  : slv116  := (others=>'1');
	constant ONES_117  : slv117  := (others=>'1'); constant ONES_118  : slv118  := (others=>'1'); constant ONES_119  : slv119  := (others=>'1'); constant ONES_120  : slv120  := (others=>'1');
	constant ONES_121  : slv121  := (others=>'1'); constant ONES_122  : slv122  := (others=>'1'); constant ONES_123  : slv123  := (others=>'1'); constant ONES_124  : slv124  := (others=>'1');
	constant ONES_125  : slv125  := (others=>'1'); constant ONES_126  : slv126  := (others=>'1'); constant ONES_127  : slv127  := (others=>'1'); constant ONES_128  : slv128  := (others=>'1');
	constant ONES_129  : slv129  := (others=>'1'); constant ONES_130  : slv130  := (others=>'1'); constant ONES_131  : slv131  := (others=>'1'); constant ONES_132  : slv132  := (others=>'1');
	constant ONES_133  : slv133  := (others=>'1'); constant ONES_134  : slv134  := (others=>'1'); constant ONES_135  : slv135  := (others=>'1'); constant ONES_136  : slv136  := (others=>'1');
	constant ONES_137  : slv137  := (others=>'1'); constant ONES_138  : slv138  := (others=>'1'); constant ONES_139  : slv139  := (others=>'1'); constant ONES_140  : slv140  := (others=>'1');
	constant ONES_141  : slv141  := (others=>'1'); constant ONES_142  : slv142  := (others=>'1'); constant ONES_143  : slv143  := (others=>'1'); constant ONES_144  : slv144  := (others=>'1');
	constant ONES_145  : slv145  := (others=>'1'); constant ONES_146  : slv146  := (others=>'1'); constant ONES_147  : slv147  := (others=>'1'); constant ONES_148  : slv148  := (others=>'1');
	constant ONES_149  : slv149  := (others=>'1'); constant ONES_150  : slv150  := (others=>'1'); constant ONES_151  : slv151  := (others=>'1'); constant ONES_152  : slv152  := (others=>'1');
	constant ONES_153  : slv153  := (others=>'1'); constant ONES_154  : slv154  := (others=>'1'); constant ONES_155  : slv155  := (others=>'1'); constant ONES_156  : slv156  := (others=>'1');
	constant ONES_157  : slv157  := (others=>'1'); constant ONES_158  : slv158  := (others=>'1'); constant ONES_159  : slv159  := (others=>'1'); constant ONES_160  : slv160  := (others=>'1');
	constant ONES_161  : slv161  := (others=>'1'); constant ONES_162  : slv162  := (others=>'1'); constant ONES_163  : slv163  := (others=>'1'); constant ONES_164  : slv164  := (others=>'1');
	constant ONES_165  : slv165  := (others=>'1'); constant ONES_166  : slv166  := (others=>'1'); constant ONES_167  : slv167  := (others=>'1'); constant ONES_168  : slv168  := (others=>'1');
	constant ONES_169  : slv169  := (others=>'1'); constant ONES_170  : slv170  := (others=>'1'); constant ONES_171  : slv171  := (others=>'1'); constant ONES_172  : slv172  := (others=>'1');
	constant ONES_173  : slv173  := (others=>'1'); constant ONES_174  : slv174  := (others=>'1'); constant ONES_175  : slv175  := (others=>'1'); constant ONES_176  : slv176  := (others=>'1');
	constant ONES_177  : slv177  := (others=>'1'); constant ONES_178  : slv178  := (others=>'1'); constant ONES_179  : slv179  := (others=>'1'); constant ONES_180  : slv180  := (others=>'1');
	constant ONES_181  : slv181  := (others=>'1'); constant ONES_182  : slv182  := (others=>'1'); constant ONES_183  : slv183  := (others=>'1'); constant ONES_184  : slv184  := (others=>'1');
	constant ONES_185  : slv185  := (others=>'1'); constant ONES_186  : slv186  := (others=>'1'); constant ONES_187  : slv187  := (others=>'1'); constant ONES_188  : slv188  := (others=>'1');
	constant ONES_189  : slv189  := (others=>'1'); constant ONES_190  : slv190  := (others=>'1'); constant ONES_191  : slv191  := (others=>'1'); constant ONES_192  : slv192  := (others=>'1');
	constant ONES_193  : slv193  := (others=>'1'); constant ONES_194  : slv194  := (others=>'1'); constant ONES_195  : slv195  := (others=>'1'); constant ONES_196  : slv196  := (others=>'1');
	constant ONES_197  : slv197  := (others=>'1'); constant ONES_198  : slv198  := (others=>'1'); constant ONES_199  : slv199  := (others=>'1'); constant ONES_200  : slv200  := (others=>'1');
	constant ONES_201  : slv201  := (others=>'1'); constant ONES_202  : slv202  := (others=>'1'); constant ONES_203  : slv203  := (others=>'1'); constant ONES_204  : slv204  := (others=>'1');
	constant ONES_205  : slv205  := (others=>'1'); constant ONES_206  : slv206  := (others=>'1'); constant ONES_207  : slv207  := (others=>'1'); constant ONES_208  : slv208  := (others=>'1');
	constant ONES_209  : slv209  := (others=>'1'); constant ONES_210  : slv210  := (others=>'1'); constant ONES_211  : slv211  := (others=>'1'); constant ONES_212  : slv212  := (others=>'1');
	constant ONES_213  : slv213  := (others=>'1'); constant ONES_214  : slv214  := (others=>'1'); constant ONES_215  : slv215  := (others=>'1'); constant ONES_216  : slv216  := (others=>'1');
	constant ONES_217  : slv217  := (others=>'1'); constant ONES_218  : slv218  := (others=>'1'); constant ONES_219  : slv219  := (others=>'1'); constant ONES_220  : slv220  := (others=>'1');
	constant ONES_221  : slv221  := (others=>'1'); constant ONES_222  : slv222  := (others=>'1'); constant ONES_223  : slv223  := (others=>'1'); constant ONES_224  : slv224  := (others=>'1');
	constant ONES_225  : slv225  := (others=>'1'); constant ONES_226  : slv226  := (others=>'1'); constant ONES_227  : slv227  := (others=>'1'); constant ONES_228  : slv228  := (others=>'1');
	constant ONES_229  : slv229  := (others=>'1'); constant ONES_230  : slv230  := (others=>'1'); constant ONES_231  : slv231  := (others=>'1'); constant ONES_232  : slv232  := (others=>'1');
	constant ONES_233  : slv233  := (others=>'1'); constant ONES_234  : slv234  := (others=>'1'); constant ONES_235  : slv235  := (others=>'1'); constant ONES_236  : slv236  := (others=>'1');
	constant ONES_237  : slv237  := (others=>'1'); constant ONES_238  : slv238  := (others=>'1'); constant ONES_239  : slv239  := (others=>'1'); constant ONES_240  : slv240  := (others=>'1');
	constant ONES_241  : slv241  := (others=>'1'); constant ONES_242  : slv242  := (others=>'1'); constant ONES_243  : slv243  := (others=>'1'); constant ONES_244  : slv244  := (others=>'1');
	constant ONES_245  : slv245  := (others=>'1'); constant ONES_246  : slv246  := (others=>'1'); constant ONES_247  : slv247  := (others=>'1'); constant ONES_248  : slv248  := (others=>'1');
	constant ONES_249  : slv249  := (others=>'1'); constant ONES_250  : slv250  := (others=>'1'); constant ONES_251  : slv251  := (others=>'1'); constant ONES_252  : slv252  := (others=>'1');
	constant ONES_253  : slv253  := (others=>'1'); constant ONES_254  : slv254  := (others=>'1'); constant ONES_255  : slv255  := (others=>'1'); constant ONES_256  : slv256  := (others=>'1');
	constant ONES_257  : slv257  := (others=>'1'); constant ONES_258  : slv258  := (others=>'1'); constant ONES_259  : slv259  := (others=>'1'); constant ONES_260  : slv260  := (others=>'1');
	constant ONES_261  : slv261  := (others=>'1'); constant ONES_262  : slv262  := (others=>'1'); constant ONES_263  : slv263  := (others=>'1'); constant ONES_264  : slv264  := (others=>'1');
	constant ONES_265  : slv265  := (others=>'1'); constant ONES_266  : slv266  := (others=>'1'); constant ONES_267  : slv267  := (others=>'1'); constant ONES_268  : slv268  := (others=>'1');
	constant ONES_269  : slv269  := (others=>'1'); constant ONES_270  : slv270  := (others=>'1'); constant ONES_271  : slv271  := (others=>'1'); constant ONES_272  : slv272  := (others=>'1');
	constant ONES_273  : slv273  := (others=>'1'); constant ONES_274  : slv274  := (others=>'1'); constant ONES_275  : slv275  := (others=>'1'); constant ONES_276  : slv276  := (others=>'1');
	constant ONES_277  : slv277  := (others=>'1'); constant ONES_278  : slv278  := (others=>'1'); constant ONES_279  : slv279  := (others=>'1'); constant ONES_280  : slv280  := (others=>'1');
	constant ONES_281  : slv281  := (others=>'1'); constant ONES_282  : slv282  := (others=>'1'); constant ONES_283  : slv283  := (others=>'1'); constant ONES_284  : slv284  := (others=>'1');
	constant ONES_285  : slv285  := (others=>'1'); constant ONES_286  : slv286  := (others=>'1'); constant ONES_287  : slv287  := (others=>'1'); constant ONES_288  : slv288  := (others=>'1');
	constant ONES_289  : slv289  := (others=>'1'); constant ONES_290  : slv290  := (others=>'1'); constant ONES_291  : slv291  := (others=>'1'); constant ONES_292  : slv292  := (others=>'1');
	constant ONES_293  : slv293  := (others=>'1'); constant ONES_294  : slv294  := (others=>'1'); constant ONES_295  : slv295  := (others=>'1'); constant ONES_296  : slv296  := (others=>'1');
	constant ONES_297  : slv297  := (others=>'1'); constant ONES_298  : slv298  := (others=>'1'); constant ONES_299  : slv299  := (others=>'1'); constant ONES_300  : slv300  := (others=>'1');
	constant ONES_301  : slv301  := (others=>'1'); constant ONES_302  : slv302  := (others=>'1'); constant ONES_303  : slv303  := (others=>'1'); constant ONES_304  : slv304  := (others=>'1');
	constant ONES_305  : slv305  := (others=>'1'); constant ONES_306  : slv306  := (others=>'1'); constant ONES_307  : slv307  := (others=>'1'); constant ONES_308  : slv308  := (others=>'1');
	constant ONES_309  : slv309  := (others=>'1'); constant ONES_310  : slv310  := (others=>'1'); constant ONES_311  : slv311  := (others=>'1'); constant ONES_312  : slv312  := (others=>'1');
	constant ONES_313  : slv313  := (others=>'1'); constant ONES_314  : slv314  := (others=>'1'); constant ONES_315  : slv315  := (others=>'1'); constant ONES_316  : slv316  := (others=>'1');
	constant ONES_317  : slv317  := (others=>'1'); constant ONES_318  : slv318  := (others=>'1'); constant ONES_319  : slv319  := (others=>'1'); constant ONES_320  : slv320  := (others=>'1');
	constant ONES_321  : slv321  := (others=>'1'); constant ONES_322  : slv322  := (others=>'1'); constant ONES_323  : slv323  := (others=>'1'); constant ONES_324  : slv324  := (others=>'1');
	constant ONES_325  : slv325  := (others=>'1'); constant ONES_326  : slv326  := (others=>'1'); constant ONES_327  : slv327  := (others=>'1'); constant ONES_328  : slv328  := (others=>'1');
	constant ONES_329  : slv329  := (others=>'1'); constant ONES_330  : slv330  := (others=>'1'); constant ONES_331  : slv331  := (others=>'1'); constant ONES_332  : slv332  := (others=>'1');
	constant ONES_333  : slv333  := (others=>'1'); constant ONES_334  : slv334  := (others=>'1'); constant ONES_335  : slv335  := (others=>'1'); constant ONES_336  : slv336  := (others=>'1');
	constant ONES_337  : slv337  := (others=>'1'); constant ONES_338  : slv338  := (others=>'1'); constant ONES_339  : slv339  := (others=>'1'); constant ONES_340  : slv340  := (others=>'1');
	constant ONES_341  : slv341  := (others=>'1'); constant ONES_342  : slv342  := (others=>'1'); constant ONES_343  : slv343  := (others=>'1'); constant ONES_344  : slv344  := (others=>'1');
	constant ONES_345  : slv345  := (others=>'1'); constant ONES_346  : slv346  := (others=>'1'); constant ONES_347  : slv347  := (others=>'1'); constant ONES_348  : slv348  := (others=>'1');
	constant ONES_349  : slv349  := (others=>'1'); constant ONES_350  : slv350  := (others=>'1'); constant ONES_351  : slv351  := (others=>'1'); constant ONES_352  : slv352  := (others=>'1');
	constant ONES_353  : slv353  := (others=>'1'); constant ONES_354  : slv354  := (others=>'1'); constant ONES_355  : slv355  := (others=>'1'); constant ONES_356  : slv356  := (others=>'1');
	constant ONES_357  : slv357  := (others=>'1'); constant ONES_358  : slv358  := (others=>'1'); constant ONES_359  : slv359  := (others=>'1'); constant ONES_360  : slv360  := (others=>'1');
	constant ONES_361  : slv361  := (others=>'1'); constant ONES_362  : slv362  := (others=>'1'); constant ONES_363  : slv363  := (others=>'1'); constant ONES_364  : slv364  := (others=>'1');
	constant ONES_365  : slv365  := (others=>'1'); constant ONES_366  : slv366  := (others=>'1'); constant ONES_367  : slv367  := (others=>'1'); constant ONES_368  : slv368  := (others=>'1');
	constant ONES_369  : slv369  := (others=>'1'); constant ONES_370  : slv370  := (others=>'1'); constant ONES_371  : slv371  := (others=>'1'); constant ONES_372  : slv372  := (others=>'1');
	constant ONES_373  : slv373  := (others=>'1'); constant ONES_374  : slv374  := (others=>'1'); constant ONES_375  : slv375  := (others=>'1'); constant ONES_376  : slv376  := (others=>'1');
	constant ONES_377  : slv377  := (others=>'1'); constant ONES_378  : slv378  := (others=>'1'); constant ONES_379  : slv379  := (others=>'1'); constant ONES_380  : slv380  := (others=>'1');
	constant ONES_381  : slv381  := (others=>'1'); constant ONES_382  : slv382  := (others=>'1'); constant ONES_383  : slv383  := (others=>'1'); constant ONES_384  : slv384  := (others=>'1');
	constant ONES_385  : slv385  := (others=>'1'); constant ONES_386  : slv386  := (others=>'1'); constant ONES_387  : slv387  := (others=>'1'); constant ONES_388  : slv388  := (others=>'1');
	constant ONES_389  : slv389  := (others=>'1'); constant ONES_390  : slv390  := (others=>'1'); constant ONES_391  : slv391  := (others=>'1'); constant ONES_392  : slv392  := (others=>'1');
	constant ONES_393  : slv393  := (others=>'1'); constant ONES_394  : slv394  := (others=>'1'); constant ONES_395  : slv395  := (others=>'1'); constant ONES_396  : slv396  := (others=>'1');
	constant ONES_397  : slv397  := (others=>'1'); constant ONES_398  : slv398  := (others=>'1'); constant ONES_399  : slv399  := (others=>'1'); constant ONES_400  : slv400  := (others=>'1');
	constant ONES_401  : slv401  := (others=>'1'); constant ONES_402  : slv402  := (others=>'1'); constant ONES_403  : slv403  := (others=>'1'); constant ONES_404  : slv404  := (others=>'1');
	constant ONES_405  : slv405  := (others=>'1'); constant ONES_406  : slv406  := (others=>'1'); constant ONES_407  : slv407  := (others=>'1'); constant ONES_408  : slv408  := (others=>'1');
	constant ONES_409  : slv409  := (others=>'1'); constant ONES_410  : slv410  := (others=>'1'); constant ONES_411  : slv411  := (others=>'1'); constant ONES_412  : slv412  := (others=>'1');
	constant ONES_413  : slv413  := (others=>'1'); constant ONES_414  : slv414  := (others=>'1'); constant ONES_415  : slv415  := (others=>'1'); constant ONES_416  : slv416  := (others=>'1');
	constant ONES_417  : slv417  := (others=>'1'); constant ONES_418  : slv418  := (others=>'1'); constant ONES_419  : slv419  := (others=>'1'); constant ONES_420  : slv420  := (others=>'1');
	constant ONES_421  : slv421  := (others=>'1'); constant ONES_422  : slv422  := (others=>'1'); constant ONES_423  : slv423  := (others=>'1'); constant ONES_424  : slv424  := (others=>'1');
	constant ONES_425  : slv425  := (others=>'1'); constant ONES_426  : slv426  := (others=>'1'); constant ONES_427  : slv427  := (others=>'1'); constant ONES_428  : slv428  := (others=>'1');
	constant ONES_429  : slv429  := (others=>'1'); constant ONES_430  : slv430  := (others=>'1'); constant ONES_431  : slv431  := (others=>'1'); constant ONES_432  : slv432  := (others=>'1');
	constant ONES_433  : slv433  := (others=>'1'); constant ONES_434  : slv434  := (others=>'1'); constant ONES_435  : slv435  := (others=>'1'); constant ONES_436  : slv436  := (others=>'1');
	constant ONES_437  : slv437  := (others=>'1'); constant ONES_438  : slv438  := (others=>'1'); constant ONES_439  : slv439  := (others=>'1'); constant ONES_440  : slv440  := (others=>'1');
	constant ONES_441  : slv441  := (others=>'1'); constant ONES_442  : slv442  := (others=>'1'); constant ONES_443  : slv443  := (others=>'1'); constant ONES_444  : slv444  := (others=>'1');
	constant ONES_445  : slv445  := (others=>'1'); constant ONES_446  : slv446  := (others=>'1'); constant ONES_447  : slv447  := (others=>'1'); constant ONES_448  : slv448  := (others=>'1');
	constant ONES_449  : slv449  := (others=>'1'); constant ONES_450  : slv450  := (others=>'1'); constant ONES_451  : slv451  := (others=>'1'); constant ONES_452  : slv452  := (others=>'1');
	constant ONES_453  : slv453  := (others=>'1'); constant ONES_454  : slv454  := (others=>'1'); constant ONES_455  : slv455  := (others=>'1'); constant ONES_456  : slv456  := (others=>'1');
	constant ONES_457  : slv457  := (others=>'1'); constant ONES_458  : slv458  := (others=>'1'); constant ONES_459  : slv459  := (others=>'1'); constant ONES_460  : slv460  := (others=>'1');
	constant ONES_461  : slv461  := (others=>'1'); constant ONES_462  : slv462  := (others=>'1'); constant ONES_463  : slv463  := (others=>'1'); constant ONES_464  : slv464  := (others=>'1');
	constant ONES_465  : slv465  := (others=>'1'); constant ONES_466  : slv466  := (others=>'1'); constant ONES_467  : slv467  := (others=>'1'); constant ONES_468  : slv468  := (others=>'1');
	constant ONES_469  : slv469  := (others=>'1'); constant ONES_470  : slv470  := (others=>'1'); constant ONES_471  : slv471  := (others=>'1'); constant ONES_472  : slv472  := (others=>'1');
	constant ONES_473  : slv473  := (others=>'1'); constant ONES_474  : slv474  := (others=>'1'); constant ONES_475  : slv475  := (others=>'1'); constant ONES_476  : slv476  := (others=>'1');
	constant ONES_477  : slv477  := (others=>'1'); constant ONES_478  : slv478  := (others=>'1'); constant ONES_479  : slv479  := (others=>'1'); constant ONES_480  : slv480  := (others=>'1');
	constant ONES_481  : slv481  := (others=>'1'); constant ONES_482  : slv482  := (others=>'1'); constant ONES_483  : slv483  := (others=>'1'); constant ONES_484  : slv484  := (others=>'1');
	constant ONES_485  : slv485  := (others=>'1'); constant ONES_486  : slv486  := (others=>'1'); constant ONES_487  : slv487  := (others=>'1'); constant ONES_488  : slv488  := (others=>'1');
	constant ONES_489  : slv489  := (others=>'1'); constant ONES_490  : slv490  := (others=>'1'); constant ONES_491  : slv491  := (others=>'1'); constant ONES_492  : slv492  := (others=>'1');
	constant ONES_493  : slv493  := (others=>'1'); constant ONES_494  : slv494  := (others=>'1'); constant ONES_495  : slv495  := (others=>'1'); constant ONES_496  : slv496  := (others=>'1');
	constant ONES_497  : slv497  := (others=>'1'); constant ONES_498  : slv498  := (others=>'1'); constant ONES_499  : slv499  := (others=>'1'); constant ONES_500  : slv500  := (others=>'1');
	constant ONES_501  : slv501  := (others=>'1'); constant ONES_502  : slv502  := (others=>'1'); constant ONES_503  : slv503  := (others=>'1'); constant ONES_504  : slv504  := (others=>'1');
	constant ONES_505  : slv505  := (others=>'1'); constant ONES_506  : slv506  := (others=>'1'); constant ONES_507  : slv507  := (others=>'1'); constant ONES_508  : slv508  := (others=>'1');
	constant ONES_509  : slv509  := (others=>'1'); constant ONES_510  : slv510  := (others=>'1'); constant ONES_511  : slv511  := (others=>'1'); constant ONES_512  : slv512  := (others=>'1');
	constant ONES_513  : slv513  := (others=>'1'); constant ONES_514  : slv514  := (others=>'1'); constant ONES_515  : slv515  := (others=>'1'); constant ONES_516  : slv516  := (others=>'1');
	constant ONES_517  : slv517  := (others=>'1'); constant ONES_518  : slv518  := (others=>'1'); constant ONES_519  : slv519  := (others=>'1'); constant ONES_520  : slv520  := (others=>'1');
	constant ONES_521  : slv521  := (others=>'1'); constant ONES_522  : slv522  := (others=>'1'); constant ONES_523  : slv523  := (others=>'1'); constant ONES_524  : slv524  := (others=>'1');
	constant ONES_525  : slv525  := (others=>'1'); constant ONES_526  : slv526  := (others=>'1'); constant ONES_527  : slv527  := (others=>'1'); constant ONES_528  : slv528  := (others=>'1');
	constant ONES_529  : slv529  := (others=>'1'); constant ONES_530  : slv530  := (others=>'1'); constant ONES_531  : slv531  := (others=>'1'); constant ONES_532  : slv532  := (others=>'1');
	constant ONES_533  : slv533  := (others=>'1'); constant ONES_534  : slv534  := (others=>'1'); constant ONES_535  : slv535  := (others=>'1'); constant ONES_536  : slv536  := (others=>'1');
	constant ONES_537  : slv537  := (others=>'1'); constant ONES_538  : slv538  := (others=>'1'); constant ONES_539  : slv539  := (others=>'1'); constant ONES_540  : slv540  := (others=>'1');
	constant ONES_541  : slv541  := (others=>'1'); constant ONES_542  : slv542  := (others=>'1'); constant ONES_543  : slv543  := (others=>'1'); constant ONES_544  : slv544  := (others=>'1');
	constant ONES_545  : slv545  := (others=>'1'); constant ONES_546  : slv546  := (others=>'1'); constant ONES_547  : slv547  := (others=>'1'); constant ONES_548  : slv548  := (others=>'1');
	constant ONES_549  : slv549  := (others=>'1'); constant ONES_550  : slv550  := (others=>'1'); constant ONES_551  : slv551  := (others=>'1'); constant ONES_552  : slv552  := (others=>'1');
	constant ONES_553  : slv553  := (others=>'1'); constant ONES_554  : slv554  := (others=>'1'); constant ONES_555  : slv555  := (others=>'1'); constant ONES_556  : slv556  := (others=>'1');
	constant ONES_557  : slv557  := (others=>'1'); constant ONES_558  : slv558  := (others=>'1'); constant ONES_559  : slv559  := (others=>'1'); constant ONES_560  : slv560  := (others=>'1');
	constant ONES_561  : slv561  := (others=>'1'); constant ONES_562  : slv562  := (others=>'1'); constant ONES_563  : slv563  := (others=>'1'); constant ONES_564  : slv564  := (others=>'1');
	constant ONES_565  : slv565  := (others=>'1'); constant ONES_566  : slv566  := (others=>'1'); constant ONES_567  : slv567  := (others=>'1'); constant ONES_568  : slv568  := (others=>'1');
	constant ONES_569  : slv569  := (others=>'1'); constant ONES_570  : slv570  := (others=>'1'); constant ONES_571  : slv571  := (others=>'1'); constant ONES_572  : slv572  := (others=>'1');
	constant ONES_573  : slv573  := (others=>'1'); constant ONES_574  : slv574  := (others=>'1'); constant ONES_575  : slv575  := (others=>'1'); constant ONES_576  : slv576  := (others=>'1');
	constant ONES_577  : slv577  := (others=>'1'); constant ONES_578  : slv578  := (others=>'1'); constant ONES_579  : slv579  := (others=>'1'); constant ONES_580  : slv580  := (others=>'1');
	constant ONES_581  : slv581  := (others=>'1'); constant ONES_582  : slv582  := (others=>'1'); constant ONES_583  : slv583  := (others=>'1'); constant ONES_584  : slv584  := (others=>'1');
	constant ONES_585  : slv585  := (others=>'1'); constant ONES_586  : slv586  := (others=>'1'); constant ONES_587  : slv587  := (others=>'1'); constant ONES_588  : slv588  := (others=>'1');
	constant ONES_589  : slv589  := (others=>'1'); constant ONES_590  : slv590  := (others=>'1'); constant ONES_591  : slv591  := (others=>'1'); constant ONES_592  : slv592  := (others=>'1');
	constant ONES_593  : slv593  := (others=>'1'); constant ONES_594  : slv594  := (others=>'1'); constant ONES_595  : slv595  := (others=>'1'); constant ONES_596  : slv596  := (others=>'1');
	constant ONES_597  : slv597  := (others=>'1'); constant ONES_598  : slv598  := (others=>'1'); constant ONES_599  : slv599  := (others=>'1'); constant ONES_600  : slv600  := (others=>'1');
	constant ONES_601  : slv601  := (others=>'1'); constant ONES_602  : slv602  := (others=>'1'); constant ONES_603  : slv603  := (others=>'1'); constant ONES_604  : slv604  := (others=>'1');
	constant ONES_605  : slv605  := (others=>'1'); constant ONES_606  : slv606  := (others=>'1'); constant ONES_607  : slv607  := (others=>'1'); constant ONES_608  : slv608  := (others=>'1');
	constant ONES_609  : slv609  := (others=>'1'); constant ONES_610  : slv610  := (others=>'1'); constant ONES_611  : slv611  := (others=>'1'); constant ONES_612  : slv612  := (others=>'1');
	constant ONES_613  : slv613  := (others=>'1'); constant ONES_614  : slv614  := (others=>'1'); constant ONES_615  : slv615  := (others=>'1'); constant ONES_616  : slv616  := (others=>'1');
	constant ONES_617  : slv617  := (others=>'1'); constant ONES_618  : slv618  := (others=>'1'); constant ONES_619  : slv619  := (others=>'1'); constant ONES_620  : slv620  := (others=>'1');
	constant ONES_621  : slv621  := (others=>'1'); constant ONES_622  : slv622  := (others=>'1'); constant ONES_623  : slv623  := (others=>'1'); constant ONES_624  : slv624  := (others=>'1');
	constant ONES_625  : slv625  := (others=>'1'); constant ONES_626  : slv626  := (others=>'1'); constant ONES_627  : slv627  := (others=>'1'); constant ONES_628  : slv628  := (others=>'1');
	constant ONES_629  : slv629  := (others=>'1'); constant ONES_630  : slv630  := (others=>'1'); constant ONES_631  : slv631  := (others=>'1'); constant ONES_632  : slv632  := (others=>'1');
	constant ONES_633  : slv633  := (others=>'1'); constant ONES_634  : slv634  := (others=>'1'); constant ONES_635  : slv635  := (others=>'1'); constant ONES_636  : slv636  := (others=>'1');
	constant ONES_637  : slv637  := (others=>'1'); constant ONES_638  : slv638  := (others=>'1'); constant ONES_639  : slv639  := (others=>'1'); constant ONES_640  : slv640  := (others=>'1');
	constant ONES_641  : slv641  := (others=>'1'); constant ONES_642  : slv642  := (others=>'1'); constant ONES_643  : slv643  := (others=>'1'); constant ONES_644  : slv644  := (others=>'1');
	constant ONES_645  : slv645  := (others=>'1'); constant ONES_646  : slv646  := (others=>'1'); constant ONES_647  : slv647  := (others=>'1'); constant ONES_648  : slv648  := (others=>'1');
	constant ONES_649  : slv649  := (others=>'1'); constant ONES_650  : slv650  := (others=>'1'); constant ONES_651  : slv651  := (others=>'1'); constant ONES_652  : slv652  := (others=>'1');
	constant ONES_653  : slv653  := (others=>'1'); constant ONES_654  : slv654  := (others=>'1'); constant ONES_655  : slv655  := (others=>'1'); constant ONES_656  : slv656  := (others=>'1');
	constant ONES_657  : slv657  := (others=>'1'); constant ONES_658  : slv658  := (others=>'1'); constant ONES_659  : slv659  := (others=>'1'); constant ONES_660  : slv660  := (others=>'1');
	constant ONES_661  : slv661  := (others=>'1'); constant ONES_662  : slv662  := (others=>'1'); constant ONES_663  : slv663  := (others=>'1'); constant ONES_664  : slv664  := (others=>'1');
	constant ONES_665  : slv665  := (others=>'1'); constant ONES_666  : slv666  := (others=>'1'); constant ONES_667  : slv667  := (others=>'1'); constant ONES_668  : slv668  := (others=>'1');
	constant ONES_669  : slv669  := (others=>'1'); constant ONES_670  : slv670  := (others=>'1'); constant ONES_671  : slv671  := (others=>'1'); constant ONES_672  : slv672  := (others=>'1');
	constant ONES_673  : slv673  := (others=>'1'); constant ONES_674  : slv674  := (others=>'1'); constant ONES_675  : slv675  := (others=>'1'); constant ONES_676  : slv676  := (others=>'1');
	constant ONES_677  : slv677  := (others=>'1'); constant ONES_678  : slv678  := (others=>'1'); constant ONES_679  : slv679  := (others=>'1'); constant ONES_680  : slv680  := (others=>'1');
	constant ONES_681  : slv681  := (others=>'1'); constant ONES_682  : slv682  := (others=>'1'); constant ONES_683  : slv683  := (others=>'1'); constant ONES_684  : slv684  := (others=>'1');
	constant ONES_685  : slv685  := (others=>'1'); constant ONES_686  : slv686  := (others=>'1'); constant ONES_687  : slv687  := (others=>'1'); constant ONES_688  : slv688  := (others=>'1');
	constant ONES_689  : slv689  := (others=>'1'); constant ONES_690  : slv690  := (others=>'1'); constant ONES_691  : slv691  := (others=>'1'); constant ONES_692  : slv692  := (others=>'1');
	constant ONES_693  : slv693  := (others=>'1'); constant ONES_694  : slv694  := (others=>'1'); constant ONES_695  : slv695  := (others=>'1'); constant ONES_696  : slv696  := (others=>'1');
	constant ONES_697  : slv697  := (others=>'1'); constant ONES_698  : slv698  := (others=>'1'); constant ONES_699  : slv699  := (others=>'1'); constant ONES_700  : slv700  := (others=>'1');
	constant ONES_701  : slv701  := (others=>'1'); constant ONES_702  : slv702  := (others=>'1'); constant ONES_703  : slv703  := (others=>'1'); constant ONES_704  : slv704  := (others=>'1');
	constant ONES_705  : slv705  := (others=>'1'); constant ONES_706  : slv706  := (others=>'1'); constant ONES_707  : slv707  := (others=>'1'); constant ONES_708  : slv708  := (others=>'1');
	constant ONES_709  : slv709  := (others=>'1'); constant ONES_710  : slv710  := (others=>'1'); constant ONES_711  : slv711  := (others=>'1'); constant ONES_712  : slv712  := (others=>'1');
	constant ONES_713  : slv713  := (others=>'1'); constant ONES_714  : slv714  := (others=>'1'); constant ONES_715  : slv715  := (others=>'1'); constant ONES_716  : slv716  := (others=>'1');
	constant ONES_717  : slv717  := (others=>'1'); constant ONES_718  : slv718  := (others=>'1'); constant ONES_719  : slv719  := (others=>'1'); constant ONES_720  : slv720  := (others=>'1');
	constant ONES_721  : slv721  := (others=>'1'); constant ONES_722  : slv722  := (others=>'1'); constant ONES_723  : slv723  := (others=>'1'); constant ONES_724  : slv724  := (others=>'1');
	constant ONES_725  : slv725  := (others=>'1'); constant ONES_726  : slv726  := (others=>'1'); constant ONES_727  : slv727  := (others=>'1'); constant ONES_728  : slv728  := (others=>'1');
	constant ONES_729  : slv729  := (others=>'1'); constant ONES_730  : slv730  := (others=>'1'); constant ONES_731  : slv731  := (others=>'1'); constant ONES_732  : slv732  := (others=>'1');
	constant ONES_733  : slv733  := (others=>'1'); constant ONES_734  : slv734  := (others=>'1'); constant ONES_735  : slv735  := (others=>'1'); constant ONES_736  : slv736  := (others=>'1');
	constant ONES_737  : slv737  := (others=>'1'); constant ONES_738  : slv738  := (others=>'1'); constant ONES_739  : slv739  := (others=>'1'); constant ONES_740  : slv740  := (others=>'1');
	constant ONES_741  : slv741  := (others=>'1'); constant ONES_742  : slv742  := (others=>'1'); constant ONES_743  : slv743  := (others=>'1'); constant ONES_744  : slv744  := (others=>'1');
	constant ONES_745  : slv745  := (others=>'1'); constant ONES_746  : slv746  := (others=>'1'); constant ONES_747  : slv747  := (others=>'1'); constant ONES_748  : slv748  := (others=>'1');
	constant ONES_749  : slv749  := (others=>'1'); constant ONES_750  : slv750  := (others=>'1'); constant ONES_751  : slv751  := (others=>'1'); constant ONES_752  : slv752  := (others=>'1');
	constant ONES_753  : slv753  := (others=>'1'); constant ONES_754  : slv754  := (others=>'1'); constant ONES_755  : slv755  := (others=>'1'); constant ONES_756  : slv756  := (others=>'1');
	constant ONES_757  : slv757  := (others=>'1'); constant ONES_758  : slv758  := (others=>'1'); constant ONES_759  : slv759  := (others=>'1'); constant ONES_760  : slv760  := (others=>'1');
	constant ONES_761  : slv761  := (others=>'1'); constant ONES_762  : slv762  := (others=>'1'); constant ONES_763  : slv763  := (others=>'1'); constant ONES_764  : slv764  := (others=>'1');
	constant ONES_765  : slv765  := (others=>'1'); constant ONES_766  : slv766  := (others=>'1'); constant ONES_767  : slv767  := (others=>'1'); constant ONES_768  : slv768  := (others=>'1');
	constant ONES_769  : slv769  := (others=>'1'); constant ONES_770  : slv770  := (others=>'1'); constant ONES_771  : slv771  := (others=>'1'); constant ONES_772  : slv772  := (others=>'1');
	constant ONES_773  : slv773  := (others=>'1'); constant ONES_774  : slv774  := (others=>'1'); constant ONES_775  : slv775  := (others=>'1'); constant ONES_776  : slv776  := (others=>'1');
	constant ONES_777  : slv777  := (others=>'1'); constant ONES_778  : slv778  := (others=>'1'); constant ONES_779  : slv779  := (others=>'1'); constant ONES_780  : slv780  := (others=>'1');
	constant ONES_781  : slv781  := (others=>'1'); constant ONES_782  : slv782  := (others=>'1'); constant ONES_783  : slv783  := (others=>'1'); constant ONES_784  : slv784  := (others=>'1');
	constant ONES_785  : slv785  := (others=>'1'); constant ONES_786  : slv786  := (others=>'1'); constant ONES_787  : slv787  := (others=>'1'); constant ONES_788  : slv788  := (others=>'1');
	constant ONES_789  : slv789  := (others=>'1'); constant ONES_790  : slv790  := (others=>'1'); constant ONES_791  : slv791  := (others=>'1'); constant ONES_792  : slv792  := (others=>'1');
	constant ONES_793  : slv793  := (others=>'1'); constant ONES_794  : slv794  := (others=>'1'); constant ONES_795  : slv795  := (others=>'1'); constant ONES_796  : slv796  := (others=>'1');
	constant ONES_797  : slv797  := (others=>'1'); constant ONES_798  : slv798  := (others=>'1'); constant ONES_799  : slv799  := (others=>'1'); constant ONES_800  : slv800  := (others=>'1');
	constant ONES_801  : slv801  := (others=>'1'); constant ONES_802  : slv802  := (others=>'1'); constant ONES_803  : slv803  := (others=>'1'); constant ONES_804  : slv804  := (others=>'1');
	constant ONES_805  : slv805  := (others=>'1'); constant ONES_806  : slv806  := (others=>'1'); constant ONES_807  : slv807  := (others=>'1'); constant ONES_808  : slv808  := (others=>'1');
	constant ONES_809  : slv809  := (others=>'1'); constant ONES_810  : slv810  := (others=>'1'); constant ONES_811  : slv811  := (others=>'1'); constant ONES_812  : slv812  := (others=>'1');
	constant ONES_813  : slv813  := (others=>'1'); constant ONES_814  : slv814  := (others=>'1'); constant ONES_815  : slv815  := (others=>'1'); constant ONES_816  : slv816  := (others=>'1');
	constant ONES_817  : slv817  := (others=>'1'); constant ONES_818  : slv818  := (others=>'1'); constant ONES_819  : slv819  := (others=>'1'); constant ONES_820  : slv820  := (others=>'1');
	constant ONES_821  : slv821  := (others=>'1'); constant ONES_822  : slv822  := (others=>'1'); constant ONES_823  : slv823  := (others=>'1'); constant ONES_824  : slv824  := (others=>'1');
	constant ONES_825  : slv825  := (others=>'1'); constant ONES_826  : slv826  := (others=>'1'); constant ONES_827  : slv827  := (others=>'1'); constant ONES_828  : slv828  := (others=>'1');
	constant ONES_829  : slv829  := (others=>'1'); constant ONES_830  : slv830  := (others=>'1'); constant ONES_831  : slv831  := (others=>'1'); constant ONES_832  : slv832  := (others=>'1');
	constant ONES_833  : slv833  := (others=>'1'); constant ONES_834  : slv834  := (others=>'1'); constant ONES_835  : slv835  := (others=>'1'); constant ONES_836  : slv836  := (others=>'1');
	constant ONES_837  : slv837  := (others=>'1'); constant ONES_838  : slv838  := (others=>'1'); constant ONES_839  : slv839  := (others=>'1'); constant ONES_840  : slv840  := (others=>'1');
	constant ONES_841  : slv841  := (others=>'1'); constant ONES_842  : slv842  := (others=>'1'); constant ONES_843  : slv843  := (others=>'1'); constant ONES_844  : slv844  := (others=>'1');
	constant ONES_845  : slv845  := (others=>'1'); constant ONES_846  : slv846  := (others=>'1'); constant ONES_847  : slv847  := (others=>'1'); constant ONES_848  : slv848  := (others=>'1');
	constant ONES_849  : slv849  := (others=>'1'); constant ONES_850  : slv850  := (others=>'1'); constant ONES_851  : slv851  := (others=>'1'); constant ONES_852  : slv852  := (others=>'1');
	constant ONES_853  : slv853  := (others=>'1'); constant ONES_854  : slv854  := (others=>'1'); constant ONES_855  : slv855  := (others=>'1'); constant ONES_856  : slv856  := (others=>'1');
	constant ONES_857  : slv857  := (others=>'1'); constant ONES_858  : slv858  := (others=>'1'); constant ONES_859  : slv859  := (others=>'1'); constant ONES_860  : slv860  := (others=>'1');
	constant ONES_861  : slv861  := (others=>'1'); constant ONES_862  : slv862  := (others=>'1'); constant ONES_863  : slv863  := (others=>'1'); constant ONES_864  : slv864  := (others=>'1');
	constant ONES_865  : slv865  := (others=>'1'); constant ONES_866  : slv866  := (others=>'1'); constant ONES_867  : slv867  := (others=>'1'); constant ONES_868  : slv868  := (others=>'1');
	constant ONES_869  : slv869  := (others=>'1'); constant ONES_870  : slv870  := (others=>'1'); constant ONES_871  : slv871  := (others=>'1'); constant ONES_872  : slv872  := (others=>'1');
	constant ONES_873  : slv873  := (others=>'1'); constant ONES_874  : slv874  := (others=>'1'); constant ONES_875  : slv875  := (others=>'1'); constant ONES_876  : slv876  := (others=>'1');
	constant ONES_877  : slv877  := (others=>'1'); constant ONES_878  : slv878  := (others=>'1'); constant ONES_879  : slv879  := (others=>'1'); constant ONES_880  : slv880  := (others=>'1');
	constant ONES_881  : slv881  := (others=>'1'); constant ONES_882  : slv882  := (others=>'1'); constant ONES_883  : slv883  := (others=>'1'); constant ONES_884  : slv884  := (others=>'1');
	constant ONES_885  : slv885  := (others=>'1'); constant ONES_886  : slv886  := (others=>'1'); constant ONES_887  : slv887  := (others=>'1'); constant ONES_888  : slv888  := (others=>'1');
	constant ONES_889  : slv889  := (others=>'1'); constant ONES_890  : slv890  := (others=>'1'); constant ONES_891  : slv891  := (others=>'1'); constant ONES_892  : slv892  := (others=>'1');
	constant ONES_893  : slv893  := (others=>'1'); constant ONES_894  : slv894  := (others=>'1'); constant ONES_895  : slv895  := (others=>'1'); constant ONES_896  : slv896  := (others=>'1');
	constant ONES_897  : slv897  := (others=>'1'); constant ONES_898  : slv898  := (others=>'1'); constant ONES_899  : slv899  := (others=>'1'); constant ONES_900  : slv900  := (others=>'1');
	constant ONES_901  : slv901  := (others=>'1'); constant ONES_902  : slv902  := (others=>'1'); constant ONES_903  : slv903  := (others=>'1'); constant ONES_904  : slv904  := (others=>'1');
	constant ONES_905  : slv905  := (others=>'1'); constant ONES_906  : slv906  := (others=>'1'); constant ONES_907  : slv907  := (others=>'1'); constant ONES_908  : slv908  := (others=>'1');
	constant ONES_909  : slv909  := (others=>'1'); constant ONES_910  : slv910  := (others=>'1'); constant ONES_911  : slv911  := (others=>'1'); constant ONES_912  : slv912  := (others=>'1');
	constant ONES_913  : slv913  := (others=>'1'); constant ONES_914  : slv914  := (others=>'1'); constant ONES_915  : slv915  := (others=>'1'); constant ONES_916  : slv916  := (others=>'1');
	constant ONES_917  : slv917  := (others=>'1'); constant ONES_918  : slv918  := (others=>'1'); constant ONES_919  : slv919  := (others=>'1'); constant ONES_920  : slv920  := (others=>'1');
	constant ONES_921  : slv921  := (others=>'1'); constant ONES_922  : slv922  := (others=>'1'); constant ONES_923  : slv923  := (others=>'1'); constant ONES_924  : slv924  := (others=>'1');
	constant ONES_925  : slv925  := (others=>'1'); constant ONES_926  : slv926  := (others=>'1'); constant ONES_927  : slv927  := (others=>'1'); constant ONES_928  : slv928  := (others=>'1');
	constant ONES_929  : slv929  := (others=>'1'); constant ONES_930  : slv930  := (others=>'1'); constant ONES_931  : slv931  := (others=>'1'); constant ONES_932  : slv932  := (others=>'1');
	constant ONES_933  : slv933  := (others=>'1'); constant ONES_934  : slv934  := (others=>'1'); constant ONES_935  : slv935  := (others=>'1'); constant ONES_936  : slv936  := (others=>'1');
	constant ONES_937  : slv937  := (others=>'1'); constant ONES_938  : slv938  := (others=>'1'); constant ONES_939  : slv939  := (others=>'1'); constant ONES_940  : slv940  := (others=>'1');
	constant ONES_941  : slv941  := (others=>'1'); constant ONES_942  : slv942  := (others=>'1'); constant ONES_943  : slv943  := (others=>'1'); constant ONES_944  : slv944  := (others=>'1');
	constant ONES_945  : slv945  := (others=>'1'); constant ONES_946  : slv946  := (others=>'1'); constant ONES_947  : slv947  := (others=>'1'); constant ONES_948  : slv948  := (others=>'1');
	constant ONES_949  : slv949  := (others=>'1'); constant ONES_950  : slv950  := (others=>'1'); constant ONES_951  : slv951  := (others=>'1'); constant ONES_952  : slv952  := (others=>'1');
	constant ONES_953  : slv953  := (others=>'1'); constant ONES_954  : slv954  := (others=>'1'); constant ONES_955  : slv955  := (others=>'1'); constant ONES_956  : slv956  := (others=>'1');
	constant ONES_957  : slv957  := (others=>'1'); constant ONES_958  : slv958  := (others=>'1'); constant ONES_959  : slv959  := (others=>'1'); constant ONES_960  : slv960  := (others=>'1');
	constant ONES_961  : slv961  := (others=>'1'); constant ONES_962  : slv962  := (others=>'1'); constant ONES_963  : slv963  := (others=>'1'); constant ONES_964  : slv964  := (others=>'1');
	constant ONES_965  : slv965  := (others=>'1'); constant ONES_966  : slv966  := (others=>'1'); constant ONES_967  : slv967  := (others=>'1'); constant ONES_968  : slv968  := (others=>'1');
	constant ONES_969  : slv969  := (others=>'1'); constant ONES_970  : slv970  := (others=>'1'); constant ONES_971  : slv971  := (others=>'1'); constant ONES_972  : slv972  := (others=>'1');
	constant ONES_973  : slv973  := (others=>'1'); constant ONES_974  : slv974  := (others=>'1'); constant ONES_975  : slv975  := (others=>'1'); constant ONES_976  : slv976  := (others=>'1');
	constant ONES_977  : slv977  := (others=>'1'); constant ONES_978  : slv978  := (others=>'1'); constant ONES_979  : slv979  := (others=>'1'); constant ONES_980  : slv980  := (others=>'1');
	constant ONES_981  : slv981  := (others=>'1'); constant ONES_982  : slv982  := (others=>'1'); constant ONES_983  : slv983  := (others=>'1'); constant ONES_984  : slv984  := (others=>'1');
	constant ONES_985  : slv985  := (others=>'1'); constant ONES_986  : slv986  := (others=>'1'); constant ONES_987  : slv987  := (others=>'1'); constant ONES_988  : slv988  := (others=>'1');
	constant ONES_989  : slv989  := (others=>'1'); constant ONES_990  : slv990  := (others=>'1'); constant ONES_991  : slv991  := (others=>'1'); constant ONES_992  : slv992  := (others=>'1');
	constant ONES_993  : slv993  := (others=>'1'); constant ONES_994  : slv994  := (others=>'1'); constant ONES_995  : slv995  := (others=>'1'); constant ONES_996  : slv996  := (others=>'1');
	constant ONES_997  : slv997  := (others=>'1'); constant ONES_998  : slv998  := (others=>'1'); constant ONES_999  : slv999  := (others=>'1'); constant ONES_1000 : slv1000 := (others=>'1');
	constant ONES_1001 : slv1001 := (others=>'1'); constant ONES_1002 : slv1002 := (others=>'1'); constant ONES_1003 : slv1003 := (others=>'1'); constant ONES_1004 : slv1004 := (others=>'1');
	constant ONES_1005 : slv1005 := (others=>'1'); constant ONES_1006 : slv1006 := (others=>'1'); constant ONES_1007 : slv1007 := (others=>'1'); constant ONES_1008 : slv1008 := (others=>'1');
	constant ONES_1009 : slv1009 := (others=>'1'); constant ONES_1010 : slv1010 := (others=>'1'); constant ONES_1011 : slv1011 := (others=>'1'); constant ONES_1012 : slv1012 := (others=>'1');
	constant ONES_1013 : slv1013 := (others=>'1'); constant ONES_1014 : slv1014 := (others=>'1'); constant ONES_1015 : slv1015 := (others=>'1'); constant ONES_1016 : slv1016 := (others=>'1');
	constant ONES_1017 : slv1017 := (others=>'1'); constant ONES_1018 : slv1018 := (others=>'1'); constant ONES_1019 : slv1019 := (others=>'1'); constant ONES_1020 : slv1020 := (others=>'1');
	constant ONES_1021 : slv1021 := (others=>'1'); constant ONES_1022 : slv1022 := (others=>'1'); constant ONES_1023 : slv1023 := (others=>'1'); constant ONES_1024 : slv1024 := (others=>'1');
--**************************************************************************************************************************************************************
-- X
--**************************************************************************************************************************************************************
	constant XS      : slv(1023 downto 0) := (others=>'X');
	constant XS_1    : slv1    := (others=>'X'); constant XS_2    : slv2    := (others=>'X'); constant XS_3    : slv3    := (others=>'X'); constant XS_4    : slv4    := (others=>'X');
	constant XS_5    : slv5    := (others=>'X'); constant XS_6    : slv6    := (others=>'X'); constant XS_7    : slv7    := (others=>'X'); constant XS_8    : slv8    := (others=>'X');
	constant XS_9    : slv9    := (others=>'X'); constant XS_10   : slv10   := (others=>'X'); constant XS_11   : slv11   := (others=>'X'); constant XS_12   : slv12   := (others=>'X');
	constant XS_13   : slv13   := (others=>'X'); constant XS_14   : slv14   := (others=>'X'); constant XS_15   : slv15   := (others=>'X'); constant XS_16   : slv16   := (others=>'X');
	constant XS_17   : slv17   := (others=>'X'); constant XS_18   : slv18   := (others=>'X'); constant XS_19   : slv19   := (others=>'X'); constant XS_20   : slv20   := (others=>'X');
	constant XS_21   : slv21   := (others=>'X'); constant XS_22   : slv22   := (others=>'X'); constant XS_23   : slv23   := (others=>'X'); constant XS_24   : slv24   := (others=>'X');
	constant XS_25   : slv25   := (others=>'X'); constant XS_26   : slv26   := (others=>'X'); constant XS_27   : slv27   := (others=>'X'); constant XS_28   : slv28   := (others=>'X');
	constant XS_29   : slv29   := (others=>'X'); constant XS_30   : slv30   := (others=>'X'); constant XS_31   : slv31   := (others=>'X'); constant XS_32   : slv32   := (others=>'X');
	constant XS_33   : slv33   := (others=>'X'); constant XS_34   : slv34   := (others=>'X'); constant XS_35   : slv35   := (others=>'X'); constant XS_36   : slv36   := (others=>'X');
	constant XS_37   : slv37   := (others=>'X'); constant XS_38   : slv38   := (others=>'X'); constant XS_39   : slv39   := (others=>'X'); constant XS_40   : slv40   := (others=>'X');
	constant XS_41   : slv41   := (others=>'X'); constant XS_42   : slv42   := (others=>'X'); constant XS_43   : slv43   := (others=>'X'); constant XS_44   : slv44   := (others=>'X');
	constant XS_45   : slv45   := (others=>'X'); constant XS_46   : slv46   := (others=>'X'); constant XS_47   : slv47   := (others=>'X'); constant XS_48   : slv48   := (others=>'X');
	constant XS_49   : slv49   := (others=>'X'); constant XS_50   : slv50   := (others=>'X'); constant XS_51   : slv51   := (others=>'X'); constant XS_52   : slv52   := (others=>'X');
	constant XS_53   : slv53   := (others=>'X'); constant XS_54   : slv54   := (others=>'X'); constant XS_55   : slv55   := (others=>'X'); constant XS_56   : slv56   := (others=>'X');
	constant XS_57   : slv57   := (others=>'X'); constant XS_58   : slv58   := (others=>'X'); constant XS_59   : slv59   := (others=>'X'); constant XS_60   : slv60   := (others=>'X');
	constant XS_61   : slv61   := (others=>'X'); constant XS_62   : slv62   := (others=>'X'); constant XS_63   : slv63   := (others=>'X'); constant XS_64   : slv64   := (others=>'X');
	constant XS_65   : slv65   := (others=>'X'); constant XS_66   : slv66   := (others=>'X'); constant XS_67   : slv67   := (others=>'X'); constant XS_68   : slv68   := (others=>'X');
	constant XS_69   : slv69   := (others=>'X'); constant XS_70   : slv70   := (others=>'X'); constant XS_71   : slv71   := (others=>'X'); constant XS_72   : slv72   := (others=>'X');
	constant XS_73   : slv73   := (others=>'X'); constant XS_74   : slv74   := (others=>'X'); constant XS_75   : slv75   := (others=>'X'); constant XS_76   : slv76   := (others=>'X');
	constant XS_77   : slv77   := (others=>'X'); constant XS_78   : slv78   := (others=>'X'); constant XS_79   : slv79   := (others=>'X'); constant XS_80   : slv80   := (others=>'X');
	constant XS_81   : slv81   := (others=>'X'); constant XS_82   : slv82   := (others=>'X'); constant XS_83   : slv83   := (others=>'X'); constant XS_84   : slv84   := (others=>'X');
	constant XS_85   : slv85   := (others=>'X'); constant XS_86   : slv86   := (others=>'X'); constant XS_87   : slv87   := (others=>'X'); constant XS_88   : slv88   := (others=>'X');
	constant XS_89   : slv89   := (others=>'X'); constant XS_90   : slv90   := (others=>'X'); constant XS_91   : slv91   := (others=>'X'); constant XS_92   : slv92   := (others=>'X');
	constant XS_93   : slv93   := (others=>'X'); constant XS_94   : slv94   := (others=>'X'); constant XS_95   : slv95   := (others=>'X'); constant XS_96   : slv96   := (others=>'X');
	constant XS_97   : slv97   := (others=>'X'); constant XS_98   : slv98   := (others=>'X'); constant XS_99   : slv99   := (others=>'X'); constant XS_100  : slv100  := (others=>'X');
	constant XS_101  : slv101  := (others=>'X'); constant XS_102  : slv102  := (others=>'X'); constant XS_103  : slv103  := (others=>'X'); constant XS_104  : slv104  := (others=>'X');
	constant XS_105  : slv105  := (others=>'X'); constant XS_106  : slv106  := (others=>'X'); constant XS_107  : slv107  := (others=>'X'); constant XS_108  : slv108  := (others=>'X');
	constant XS_109  : slv109  := (others=>'X'); constant XS_110  : slv110  := (others=>'X'); constant XS_111  : slv111  := (others=>'X'); constant XS_112  : slv112  := (others=>'X');
	constant XS_113  : slv113  := (others=>'X'); constant XS_114  : slv114  := (others=>'X'); constant XS_115  : slv115  := (others=>'X'); constant XS_116  : slv116  := (others=>'X');
	constant XS_117  : slv117  := (others=>'X'); constant XS_118  : slv118  := (others=>'X'); constant XS_119  : slv119  := (others=>'X'); constant XS_120  : slv120  := (others=>'X');
	constant XS_121  : slv121  := (others=>'X'); constant XS_122  : slv122  := (others=>'X'); constant XS_123  : slv123  := (others=>'X'); constant XS_124  : slv124  := (others=>'X');
	constant XS_125  : slv125  := (others=>'X'); constant XS_126  : slv126  := (others=>'X'); constant XS_127  : slv127  := (others=>'X'); constant XS_128  : slv128  := (others=>'X');
	constant XS_129  : slv129  := (others=>'X'); constant XS_130  : slv130  := (others=>'X'); constant XS_131  : slv131  := (others=>'X'); constant XS_132  : slv132  := (others=>'X');
	constant XS_133  : slv133  := (others=>'X'); constant XS_134  : slv134  := (others=>'X'); constant XS_135  : slv135  := (others=>'X'); constant XS_136  : slv136  := (others=>'X');
	constant XS_137  : slv137  := (others=>'X'); constant XS_138  : slv138  := (others=>'X'); constant XS_139  : slv139  := (others=>'X'); constant XS_140  : slv140  := (others=>'X');
	constant XS_141  : slv141  := (others=>'X'); constant XS_142  : slv142  := (others=>'X'); constant XS_143  : slv143  := (others=>'X'); constant XS_144  : slv144  := (others=>'X');
	constant XS_145  : slv145  := (others=>'X'); constant XS_146  : slv146  := (others=>'X'); constant XS_147  : slv147  := (others=>'X'); constant XS_148  : slv148  := (others=>'X');
	constant XS_149  : slv149  := (others=>'X'); constant XS_150  : slv150  := (others=>'X'); constant XS_151  : slv151  := (others=>'X'); constant XS_152  : slv152  := (others=>'X');
	constant XS_153  : slv153  := (others=>'X'); constant XS_154  : slv154  := (others=>'X'); constant XS_155  : slv155  := (others=>'X'); constant XS_156  : slv156  := (others=>'X');
	constant XS_157  : slv157  := (others=>'X'); constant XS_158  : slv158  := (others=>'X'); constant XS_159  : slv159  := (others=>'X'); constant XS_160  : slv160  := (others=>'X');
	constant XS_161  : slv161  := (others=>'X'); constant XS_162  : slv162  := (others=>'X'); constant XS_163  : slv163  := (others=>'X'); constant XS_164  : slv164  := (others=>'X');
	constant XS_165  : slv165  := (others=>'X'); constant XS_166  : slv166  := (others=>'X'); constant XS_167  : slv167  := (others=>'X'); constant XS_168  : slv168  := (others=>'X');
	constant XS_169  : slv169  := (others=>'X'); constant XS_170  : slv170  := (others=>'X'); constant XS_171  : slv171  := (others=>'X'); constant XS_172  : slv172  := (others=>'X');
	constant XS_173  : slv173  := (others=>'X'); constant XS_174  : slv174  := (others=>'X'); constant XS_175  : slv175  := (others=>'X'); constant XS_176  : slv176  := (others=>'X');
	constant XS_177  : slv177  := (others=>'X'); constant XS_178  : slv178  := (others=>'X'); constant XS_179  : slv179  := (others=>'X'); constant XS_180  : slv180  := (others=>'X');
	constant XS_181  : slv181  := (others=>'X'); constant XS_182  : slv182  := (others=>'X'); constant XS_183  : slv183  := (others=>'X'); constant XS_184  : slv184  := (others=>'X');
	constant XS_185  : slv185  := (others=>'X'); constant XS_186  : slv186  := (others=>'X'); constant XS_187  : slv187  := (others=>'X'); constant XS_188  : slv188  := (others=>'X');
	constant XS_189  : slv189  := (others=>'X'); constant XS_190  : slv190  := (others=>'X'); constant XS_191  : slv191  := (others=>'X'); constant XS_192  : slv192  := (others=>'X');
	constant XS_193  : slv193  := (others=>'X'); constant XS_194  : slv194  := (others=>'X'); constant XS_195  : slv195  := (others=>'X'); constant XS_196  : slv196  := (others=>'X');
	constant XS_197  : slv197  := (others=>'X'); constant XS_198  : slv198  := (others=>'X'); constant XS_199  : slv199  := (others=>'X'); constant XS_200  : slv200  := (others=>'X');
	constant XS_201  : slv201  := (others=>'X'); constant XS_202  : slv202  := (others=>'X'); constant XS_203  : slv203  := (others=>'X'); constant XS_204  : slv204  := (others=>'X');
	constant XS_205  : slv205  := (others=>'X'); constant XS_206  : slv206  := (others=>'X'); constant XS_207  : slv207  := (others=>'X'); constant XS_208  : slv208  := (others=>'X');
	constant XS_209  : slv209  := (others=>'X'); constant XS_210  : slv210  := (others=>'X'); constant XS_211  : slv211  := (others=>'X'); constant XS_212  : slv212  := (others=>'X');
	constant XS_213  : slv213  := (others=>'X'); constant XS_214  : slv214  := (others=>'X'); constant XS_215  : slv215  := (others=>'X'); constant XS_216  : slv216  := (others=>'X');
	constant XS_217  : slv217  := (others=>'X'); constant XS_218  : slv218  := (others=>'X'); constant XS_219  : slv219  := (others=>'X'); constant XS_220  : slv220  := (others=>'X');
	constant XS_221  : slv221  := (others=>'X'); constant XS_222  : slv222  := (others=>'X'); constant XS_223  : slv223  := (others=>'X'); constant XS_224  : slv224  := (others=>'X');
	constant XS_225  : slv225  := (others=>'X'); constant XS_226  : slv226  := (others=>'X'); constant XS_227  : slv227  := (others=>'X'); constant XS_228  : slv228  := (others=>'X');
	constant XS_229  : slv229  := (others=>'X'); constant XS_230  : slv230  := (others=>'X'); constant XS_231  : slv231  := (others=>'X'); constant XS_232  : slv232  := (others=>'X');
	constant XS_233  : slv233  := (others=>'X'); constant XS_234  : slv234  := (others=>'X'); constant XS_235  : slv235  := (others=>'X'); constant XS_236  : slv236  := (others=>'X');
	constant XS_237  : slv237  := (others=>'X'); constant XS_238  : slv238  := (others=>'X'); constant XS_239  : slv239  := (others=>'X'); constant XS_240  : slv240  := (others=>'X');
	constant XS_241  : slv241  := (others=>'X'); constant XS_242  : slv242  := (others=>'X'); constant XS_243  : slv243  := (others=>'X'); constant XS_244  : slv244  := (others=>'X');
	constant XS_245  : slv245  := (others=>'X'); constant XS_246  : slv246  := (others=>'X'); constant XS_247  : slv247  := (others=>'X'); constant XS_248  : slv248  := (others=>'X');
	constant XS_249  : slv249  := (others=>'X'); constant XS_250  : slv250  := (others=>'X'); constant XS_251  : slv251  := (others=>'X'); constant XS_252  : slv252  := (others=>'X');
	constant XS_253  : slv253  := (others=>'X'); constant XS_254  : slv254  := (others=>'X'); constant XS_255  : slv255  := (others=>'X'); constant XS_256  : slv256  := (others=>'X');
	constant XS_257  : slv257  := (others=>'X'); constant XS_258  : slv258  := (others=>'X'); constant XS_259  : slv259  := (others=>'X'); constant XS_260  : slv260  := (others=>'X');
	constant XS_261  : slv261  := (others=>'X'); constant XS_262  : slv262  := (others=>'X'); constant XS_263  : slv263  := (others=>'X'); constant XS_264  : slv264  := (others=>'X');
	constant XS_265  : slv265  := (others=>'X'); constant XS_266  : slv266  := (others=>'X'); constant XS_267  : slv267  := (others=>'X'); constant XS_268  : slv268  := (others=>'X');
	constant XS_269  : slv269  := (others=>'X'); constant XS_270  : slv270  := (others=>'X'); constant XS_271  : slv271  := (others=>'X'); constant XS_272  : slv272  := (others=>'X');
	constant XS_273  : slv273  := (others=>'X'); constant XS_274  : slv274  := (others=>'X'); constant XS_275  : slv275  := (others=>'X'); constant XS_276  : slv276  := (others=>'X');
	constant XS_277  : slv277  := (others=>'X'); constant XS_278  : slv278  := (others=>'X'); constant XS_279  : slv279  := (others=>'X'); constant XS_280  : slv280  := (others=>'X');
	constant XS_281  : slv281  := (others=>'X'); constant XS_282  : slv282  := (others=>'X'); constant XS_283  : slv283  := (others=>'X'); constant XS_284  : slv284  := (others=>'X');
	constant XS_285  : slv285  := (others=>'X'); constant XS_286  : slv286  := (others=>'X'); constant XS_287  : slv287  := (others=>'X'); constant XS_288  : slv288  := (others=>'X');
	constant XS_289  : slv289  := (others=>'X'); constant XS_290  : slv290  := (others=>'X'); constant XS_291  : slv291  := (others=>'X'); constant XS_292  : slv292  := (others=>'X');
	constant XS_293  : slv293  := (others=>'X'); constant XS_294  : slv294  := (others=>'X'); constant XS_295  : slv295  := (others=>'X'); constant XS_296  : slv296  := (others=>'X');
	constant XS_297  : slv297  := (others=>'X'); constant XS_298  : slv298  := (others=>'X'); constant XS_299  : slv299  := (others=>'X'); constant XS_300  : slv300  := (others=>'X');
	constant XS_301  : slv301  := (others=>'X'); constant XS_302  : slv302  := (others=>'X'); constant XS_303  : slv303  := (others=>'X'); constant XS_304  : slv304  := (others=>'X');
	constant XS_305  : slv305  := (others=>'X'); constant XS_306  : slv306  := (others=>'X'); constant XS_307  : slv307  := (others=>'X'); constant XS_308  : slv308  := (others=>'X');
	constant XS_309  : slv309  := (others=>'X'); constant XS_310  : slv310  := (others=>'X'); constant XS_311  : slv311  := (others=>'X'); constant XS_312  : slv312  := (others=>'X');
	constant XS_313  : slv313  := (others=>'X'); constant XS_314  : slv314  := (others=>'X'); constant XS_315  : slv315  := (others=>'X'); constant XS_316  : slv316  := (others=>'X');
	constant XS_317  : slv317  := (others=>'X'); constant XS_318  : slv318  := (others=>'X'); constant XS_319  : slv319  := (others=>'X'); constant XS_320  : slv320  := (others=>'X');
	constant XS_321  : slv321  := (others=>'X'); constant XS_322  : slv322  := (others=>'X'); constant XS_323  : slv323  := (others=>'X'); constant XS_324  : slv324  := (others=>'X');
	constant XS_325  : slv325  := (others=>'X'); constant XS_326  : slv326  := (others=>'X'); constant XS_327  : slv327  := (others=>'X'); constant XS_328  : slv328  := (others=>'X');
	constant XS_329  : slv329  := (others=>'X'); constant XS_330  : slv330  := (others=>'X'); constant XS_331  : slv331  := (others=>'X'); constant XS_332  : slv332  := (others=>'X');
	constant XS_333  : slv333  := (others=>'X'); constant XS_334  : slv334  := (others=>'X'); constant XS_335  : slv335  := (others=>'X'); constant XS_336  : slv336  := (others=>'X');
	constant XS_337  : slv337  := (others=>'X'); constant XS_338  : slv338  := (others=>'X'); constant XS_339  : slv339  := (others=>'X'); constant XS_340  : slv340  := (others=>'X');
	constant XS_341  : slv341  := (others=>'X'); constant XS_342  : slv342  := (others=>'X'); constant XS_343  : slv343  := (others=>'X'); constant XS_344  : slv344  := (others=>'X');
	constant XS_345  : slv345  := (others=>'X'); constant XS_346  : slv346  := (others=>'X'); constant XS_347  : slv347  := (others=>'X'); constant XS_348  : slv348  := (others=>'X');
	constant XS_349  : slv349  := (others=>'X'); constant XS_350  : slv350  := (others=>'X'); constant XS_351  : slv351  := (others=>'X'); constant XS_352  : slv352  := (others=>'X');
	constant XS_353  : slv353  := (others=>'X'); constant XS_354  : slv354  := (others=>'X'); constant XS_355  : slv355  := (others=>'X'); constant XS_356  : slv356  := (others=>'X');
	constant XS_357  : slv357  := (others=>'X'); constant XS_358  : slv358  := (others=>'X'); constant XS_359  : slv359  := (others=>'X'); constant XS_360  : slv360  := (others=>'X');
	constant XS_361  : slv361  := (others=>'X'); constant XS_362  : slv362  := (others=>'X'); constant XS_363  : slv363  := (others=>'X'); constant XS_364  : slv364  := (others=>'X');
	constant XS_365  : slv365  := (others=>'X'); constant XS_366  : slv366  := (others=>'X'); constant XS_367  : slv367  := (others=>'X'); constant XS_368  : slv368  := (others=>'X');
	constant XS_369  : slv369  := (others=>'X'); constant XS_370  : slv370  := (others=>'X'); constant XS_371  : slv371  := (others=>'X'); constant XS_372  : slv372  := (others=>'X');
	constant XS_373  : slv373  := (others=>'X'); constant XS_374  : slv374  := (others=>'X'); constant XS_375  : slv375  := (others=>'X'); constant XS_376  : slv376  := (others=>'X');
	constant XS_377  : slv377  := (others=>'X'); constant XS_378  : slv378  := (others=>'X'); constant XS_379  : slv379  := (others=>'X'); constant XS_380  : slv380  := (others=>'X');
	constant XS_381  : slv381  := (others=>'X'); constant XS_382  : slv382  := (others=>'X'); constant XS_383  : slv383  := (others=>'X'); constant XS_384  : slv384  := (others=>'X');
	constant XS_385  : slv385  := (others=>'X'); constant XS_386  : slv386  := (others=>'X'); constant XS_387  : slv387  := (others=>'X'); constant XS_388  : slv388  := (others=>'X');
	constant XS_389  : slv389  := (others=>'X'); constant XS_390  : slv390  := (others=>'X'); constant XS_391  : slv391  := (others=>'X'); constant XS_392  : slv392  := (others=>'X');
	constant XS_393  : slv393  := (others=>'X'); constant XS_394  : slv394  := (others=>'X'); constant XS_395  : slv395  := (others=>'X'); constant XS_396  : slv396  := (others=>'X');
	constant XS_397  : slv397  := (others=>'X'); constant XS_398  : slv398  := (others=>'X'); constant XS_399  : slv399  := (others=>'X'); constant XS_400  : slv400  := (others=>'X');
	constant XS_401  : slv401  := (others=>'X'); constant XS_402  : slv402  := (others=>'X'); constant XS_403  : slv403  := (others=>'X'); constant XS_404  : slv404  := (others=>'X');
	constant XS_405  : slv405  := (others=>'X'); constant XS_406  : slv406  := (others=>'X'); constant XS_407  : slv407  := (others=>'X'); constant XS_408  : slv408  := (others=>'X');
	constant XS_409  : slv409  := (others=>'X'); constant XS_410  : slv410  := (others=>'X'); constant XS_411  : slv411  := (others=>'X'); constant XS_412  : slv412  := (others=>'X');
	constant XS_413  : slv413  := (others=>'X'); constant XS_414  : slv414  := (others=>'X'); constant XS_415  : slv415  := (others=>'X'); constant XS_416  : slv416  := (others=>'X');
	constant XS_417  : slv417  := (others=>'X'); constant XS_418  : slv418  := (others=>'X'); constant XS_419  : slv419  := (others=>'X'); constant XS_420  : slv420  := (others=>'X');
	constant XS_421  : slv421  := (others=>'X'); constant XS_422  : slv422  := (others=>'X'); constant XS_423  : slv423  := (others=>'X'); constant XS_424  : slv424  := (others=>'X');
	constant XS_425  : slv425  := (others=>'X'); constant XS_426  : slv426  := (others=>'X'); constant XS_427  : slv427  := (others=>'X'); constant XS_428  : slv428  := (others=>'X');
	constant XS_429  : slv429  := (others=>'X'); constant XS_430  : slv430  := (others=>'X'); constant XS_431  : slv431  := (others=>'X'); constant XS_432  : slv432  := (others=>'X');
	constant XS_433  : slv433  := (others=>'X'); constant XS_434  : slv434  := (others=>'X'); constant XS_435  : slv435  := (others=>'X'); constant XS_436  : slv436  := (others=>'X');
	constant XS_437  : slv437  := (others=>'X'); constant XS_438  : slv438  := (others=>'X'); constant XS_439  : slv439  := (others=>'X'); constant XS_440  : slv440  := (others=>'X');
	constant XS_441  : slv441  := (others=>'X'); constant XS_442  : slv442  := (others=>'X'); constant XS_443  : slv443  := (others=>'X'); constant XS_444  : slv444  := (others=>'X');
	constant XS_445  : slv445  := (others=>'X'); constant XS_446  : slv446  := (others=>'X'); constant XS_447  : slv447  := (others=>'X'); constant XS_448  : slv448  := (others=>'X');
	constant XS_449  : slv449  := (others=>'X'); constant XS_450  : slv450  := (others=>'X'); constant XS_451  : slv451  := (others=>'X'); constant XS_452  : slv452  := (others=>'X');
	constant XS_453  : slv453  := (others=>'X'); constant XS_454  : slv454  := (others=>'X'); constant XS_455  : slv455  := (others=>'X'); constant XS_456  : slv456  := (others=>'X');
	constant XS_457  : slv457  := (others=>'X'); constant XS_458  : slv458  := (others=>'X'); constant XS_459  : slv459  := (others=>'X'); constant XS_460  : slv460  := (others=>'X');
	constant XS_461  : slv461  := (others=>'X'); constant XS_462  : slv462  := (others=>'X'); constant XS_463  : slv463  := (others=>'X'); constant XS_464  : slv464  := (others=>'X');
	constant XS_465  : slv465  := (others=>'X'); constant XS_466  : slv466  := (others=>'X'); constant XS_467  : slv467  := (others=>'X'); constant XS_468  : slv468  := (others=>'X');
	constant XS_469  : slv469  := (others=>'X'); constant XS_470  : slv470  := (others=>'X'); constant XS_471  : slv471  := (others=>'X'); constant XS_472  : slv472  := (others=>'X');
	constant XS_473  : slv473  := (others=>'X'); constant XS_474  : slv474  := (others=>'X'); constant XS_475  : slv475  := (others=>'X'); constant XS_476  : slv476  := (others=>'X');
	constant XS_477  : slv477  := (others=>'X'); constant XS_478  : slv478  := (others=>'X'); constant XS_479  : slv479  := (others=>'X'); constant XS_480  : slv480  := (others=>'X');
	constant XS_481  : slv481  := (others=>'X'); constant XS_482  : slv482  := (others=>'X'); constant XS_483  : slv483  := (others=>'X'); constant XS_484  : slv484  := (others=>'X');
	constant XS_485  : slv485  := (others=>'X'); constant XS_486  : slv486  := (others=>'X'); constant XS_487  : slv487  := (others=>'X'); constant XS_488  : slv488  := (others=>'X');
	constant XS_489  : slv489  := (others=>'X'); constant XS_490  : slv490  := (others=>'X'); constant XS_491  : slv491  := (others=>'X'); constant XS_492  : slv492  := (others=>'X');
	constant XS_493  : slv493  := (others=>'X'); constant XS_494  : slv494  := (others=>'X'); constant XS_495  : slv495  := (others=>'X'); constant XS_496  : slv496  := (others=>'X');
	constant XS_497  : slv497  := (others=>'X'); constant XS_498  : slv498  := (others=>'X'); constant XS_499  : slv499  := (others=>'X'); constant XS_500  : slv500  := (others=>'X');
	constant XS_501  : slv501  := (others=>'X'); constant XS_502  : slv502  := (others=>'X'); constant XS_503  : slv503  := (others=>'X'); constant XS_504  : slv504  := (others=>'X');
	constant XS_505  : slv505  := (others=>'X'); constant XS_506  : slv506  := (others=>'X'); constant XS_507  : slv507  := (others=>'X'); constant XS_508  : slv508  := (others=>'X');
	constant XS_509  : slv509  := (others=>'X'); constant XS_510  : slv510  := (others=>'X'); constant XS_511  : slv511  := (others=>'X'); constant XS_512  : slv512  := (others=>'X');
	constant XS_513  : slv513  := (others=>'X'); constant XS_514  : slv514  := (others=>'X'); constant XS_515  : slv515  := (others=>'X'); constant XS_516  : slv516  := (others=>'X');
	constant XS_517  : slv517  := (others=>'X'); constant XS_518  : slv518  := (others=>'X'); constant XS_519  : slv519  := (others=>'X'); constant XS_520  : slv520  := (others=>'X');
	constant XS_521  : slv521  := (others=>'X'); constant XS_522  : slv522  := (others=>'X'); constant XS_523  : slv523  := (others=>'X'); constant XS_524  : slv524  := (others=>'X');
	constant XS_525  : slv525  := (others=>'X'); constant XS_526  : slv526  := (others=>'X'); constant XS_527  : slv527  := (others=>'X'); constant XS_528  : slv528  := (others=>'X');
	constant XS_529  : slv529  := (others=>'X'); constant XS_530  : slv530  := (others=>'X'); constant XS_531  : slv531  := (others=>'X'); constant XS_532  : slv532  := (others=>'X');
	constant XS_533  : slv533  := (others=>'X'); constant XS_534  : slv534  := (others=>'X'); constant XS_535  : slv535  := (others=>'X'); constant XS_536  : slv536  := (others=>'X');
	constant XS_537  : slv537  := (others=>'X'); constant XS_538  : slv538  := (others=>'X'); constant XS_539  : slv539  := (others=>'X'); constant XS_540  : slv540  := (others=>'X');
	constant XS_541  : slv541  := (others=>'X'); constant XS_542  : slv542  := (others=>'X'); constant XS_543  : slv543  := (others=>'X'); constant XS_544  : slv544  := (others=>'X');
	constant XS_545  : slv545  := (others=>'X'); constant XS_546  : slv546  := (others=>'X'); constant XS_547  : slv547  := (others=>'X'); constant XS_548  : slv548  := (others=>'X');
	constant XS_549  : slv549  := (others=>'X'); constant XS_550  : slv550  := (others=>'X'); constant XS_551  : slv551  := (others=>'X'); constant XS_552  : slv552  := (others=>'X');
	constant XS_553  : slv553  := (others=>'X'); constant XS_554  : slv554  := (others=>'X'); constant XS_555  : slv555  := (others=>'X'); constant XS_556  : slv556  := (others=>'X');
	constant XS_557  : slv557  := (others=>'X'); constant XS_558  : slv558  := (others=>'X'); constant XS_559  : slv559  := (others=>'X'); constant XS_560  : slv560  := (others=>'X');
	constant XS_561  : slv561  := (others=>'X'); constant XS_562  : slv562  := (others=>'X'); constant XS_563  : slv563  := (others=>'X'); constant XS_564  : slv564  := (others=>'X');
	constant XS_565  : slv565  := (others=>'X'); constant XS_566  : slv566  := (others=>'X'); constant XS_567  : slv567  := (others=>'X'); constant XS_568  : slv568  := (others=>'X');
	constant XS_569  : slv569  := (others=>'X'); constant XS_570  : slv570  := (others=>'X'); constant XS_571  : slv571  := (others=>'X'); constant XS_572  : slv572  := (others=>'X');
	constant XS_573  : slv573  := (others=>'X'); constant XS_574  : slv574  := (others=>'X'); constant XS_575  : slv575  := (others=>'X'); constant XS_576  : slv576  := (others=>'X');
	constant XS_577  : slv577  := (others=>'X'); constant XS_578  : slv578  := (others=>'X'); constant XS_579  : slv579  := (others=>'X'); constant XS_580  : slv580  := (others=>'X');
	constant XS_581  : slv581  := (others=>'X'); constant XS_582  : slv582  := (others=>'X'); constant XS_583  : slv583  := (others=>'X'); constant XS_584  : slv584  := (others=>'X');
	constant XS_585  : slv585  := (others=>'X'); constant XS_586  : slv586  := (others=>'X'); constant XS_587  : slv587  := (others=>'X'); constant XS_588  : slv588  := (others=>'X');
	constant XS_589  : slv589  := (others=>'X'); constant XS_590  : slv590  := (others=>'X'); constant XS_591  : slv591  := (others=>'X'); constant XS_592  : slv592  := (others=>'X');
	constant XS_593  : slv593  := (others=>'X'); constant XS_594  : slv594  := (others=>'X'); constant XS_595  : slv595  := (others=>'X'); constant XS_596  : slv596  := (others=>'X');
	constant XS_597  : slv597  := (others=>'X'); constant XS_598  : slv598  := (others=>'X'); constant XS_599  : slv599  := (others=>'X'); constant XS_600  : slv600  := (others=>'X');
	constant XS_601  : slv601  := (others=>'X'); constant XS_602  : slv602  := (others=>'X'); constant XS_603  : slv603  := (others=>'X'); constant XS_604  : slv604  := (others=>'X');
	constant XS_605  : slv605  := (others=>'X'); constant XS_606  : slv606  := (others=>'X'); constant XS_607  : slv607  := (others=>'X'); constant XS_608  : slv608  := (others=>'X');
	constant XS_609  : slv609  := (others=>'X'); constant XS_610  : slv610  := (others=>'X'); constant XS_611  : slv611  := (others=>'X'); constant XS_612  : slv612  := (others=>'X');
	constant XS_613  : slv613  := (others=>'X'); constant XS_614  : slv614  := (others=>'X'); constant XS_615  : slv615  := (others=>'X'); constant XS_616  : slv616  := (others=>'X');
	constant XS_617  : slv617  := (others=>'X'); constant XS_618  : slv618  := (others=>'X'); constant XS_619  : slv619  := (others=>'X'); constant XS_620  : slv620  := (others=>'X');
	constant XS_621  : slv621  := (others=>'X'); constant XS_622  : slv622  := (others=>'X'); constant XS_623  : slv623  := (others=>'X'); constant XS_624  : slv624  := (others=>'X');
	constant XS_625  : slv625  := (others=>'X'); constant XS_626  : slv626  := (others=>'X'); constant XS_627  : slv627  := (others=>'X'); constant XS_628  : slv628  := (others=>'X');
	constant XS_629  : slv629  := (others=>'X'); constant XS_630  : slv630  := (others=>'X'); constant XS_631  : slv631  := (others=>'X'); constant XS_632  : slv632  := (others=>'X');
	constant XS_633  : slv633  := (others=>'X'); constant XS_634  : slv634  := (others=>'X'); constant XS_635  : slv635  := (others=>'X'); constant XS_636  : slv636  := (others=>'X');
	constant XS_637  : slv637  := (others=>'X'); constant XS_638  : slv638  := (others=>'X'); constant XS_639  : slv639  := (others=>'X'); constant XS_640  : slv640  := (others=>'X');
	constant XS_641  : slv641  := (others=>'X'); constant XS_642  : slv642  := (others=>'X'); constant XS_643  : slv643  := (others=>'X'); constant XS_644  : slv644  := (others=>'X');
	constant XS_645  : slv645  := (others=>'X'); constant XS_646  : slv646  := (others=>'X'); constant XS_647  : slv647  := (others=>'X'); constant XS_648  : slv648  := (others=>'X');
	constant XS_649  : slv649  := (others=>'X'); constant XS_650  : slv650  := (others=>'X'); constant XS_651  : slv651  := (others=>'X'); constant XS_652  : slv652  := (others=>'X');
	constant XS_653  : slv653  := (others=>'X'); constant XS_654  : slv654  := (others=>'X'); constant XS_655  : slv655  := (others=>'X'); constant XS_656  : slv656  := (others=>'X');
	constant XS_657  : slv657  := (others=>'X'); constant XS_658  : slv658  := (others=>'X'); constant XS_659  : slv659  := (others=>'X'); constant XS_660  : slv660  := (others=>'X');
	constant XS_661  : slv661  := (others=>'X'); constant XS_662  : slv662  := (others=>'X'); constant XS_663  : slv663  := (others=>'X'); constant XS_664  : slv664  := (others=>'X');
	constant XS_665  : slv665  := (others=>'X'); constant XS_666  : slv666  := (others=>'X'); constant XS_667  : slv667  := (others=>'X'); constant XS_668  : slv668  := (others=>'X');
	constant XS_669  : slv669  := (others=>'X'); constant XS_670  : slv670  := (others=>'X'); constant XS_671  : slv671  := (others=>'X'); constant XS_672  : slv672  := (others=>'X');
	constant XS_673  : slv673  := (others=>'X'); constant XS_674  : slv674  := (others=>'X'); constant XS_675  : slv675  := (others=>'X'); constant XS_676  : slv676  := (others=>'X');
	constant XS_677  : slv677  := (others=>'X'); constant XS_678  : slv678  := (others=>'X'); constant XS_679  : slv679  := (others=>'X'); constant XS_680  : slv680  := (others=>'X');
	constant XS_681  : slv681  := (others=>'X'); constant XS_682  : slv682  := (others=>'X'); constant XS_683  : slv683  := (others=>'X'); constant XS_684  : slv684  := (others=>'X');
	constant XS_685  : slv685  := (others=>'X'); constant XS_686  : slv686  := (others=>'X'); constant XS_687  : slv687  := (others=>'X'); constant XS_688  : slv688  := (others=>'X');
	constant XS_689  : slv689  := (others=>'X'); constant XS_690  : slv690  := (others=>'X'); constant XS_691  : slv691  := (others=>'X'); constant XS_692  : slv692  := (others=>'X');
	constant XS_693  : slv693  := (others=>'X'); constant XS_694  : slv694  := (others=>'X'); constant XS_695  : slv695  := (others=>'X'); constant XS_696  : slv696  := (others=>'X');
	constant XS_697  : slv697  := (others=>'X'); constant XS_698  : slv698  := (others=>'X'); constant XS_699  : slv699  := (others=>'X'); constant XS_700  : slv700  := (others=>'X');
	constant XS_701  : slv701  := (others=>'X'); constant XS_702  : slv702  := (others=>'X'); constant XS_703  : slv703  := (others=>'X'); constant XS_704  : slv704  := (others=>'X');
	constant XS_705  : slv705  := (others=>'X'); constant XS_706  : slv706  := (others=>'X'); constant XS_707  : slv707  := (others=>'X'); constant XS_708  : slv708  := (others=>'X');
	constant XS_709  : slv709  := (others=>'X'); constant XS_710  : slv710  := (others=>'X'); constant XS_711  : slv711  := (others=>'X'); constant XS_712  : slv712  := (others=>'X');
	constant XS_713  : slv713  := (others=>'X'); constant XS_714  : slv714  := (others=>'X'); constant XS_715  : slv715  := (others=>'X'); constant XS_716  : slv716  := (others=>'X');
	constant XS_717  : slv717  := (others=>'X'); constant XS_718  : slv718  := (others=>'X'); constant XS_719  : slv719  := (others=>'X'); constant XS_720  : slv720  := (others=>'X');
	constant XS_721  : slv721  := (others=>'X'); constant XS_722  : slv722  := (others=>'X'); constant XS_723  : slv723  := (others=>'X'); constant XS_724  : slv724  := (others=>'X');
	constant XS_725  : slv725  := (others=>'X'); constant XS_726  : slv726  := (others=>'X'); constant XS_727  : slv727  := (others=>'X'); constant XS_728  : slv728  := (others=>'X');
	constant XS_729  : slv729  := (others=>'X'); constant XS_730  : slv730  := (others=>'X'); constant XS_731  : slv731  := (others=>'X'); constant XS_732  : slv732  := (others=>'X');
	constant XS_733  : slv733  := (others=>'X'); constant XS_734  : slv734  := (others=>'X'); constant XS_735  : slv735  := (others=>'X'); constant XS_736  : slv736  := (others=>'X');
	constant XS_737  : slv737  := (others=>'X'); constant XS_738  : slv738  := (others=>'X'); constant XS_739  : slv739  := (others=>'X'); constant XS_740  : slv740  := (others=>'X');
	constant XS_741  : slv741  := (others=>'X'); constant XS_742  : slv742  := (others=>'X'); constant XS_743  : slv743  := (others=>'X'); constant XS_744  : slv744  := (others=>'X');
	constant XS_745  : slv745  := (others=>'X'); constant XS_746  : slv746  := (others=>'X'); constant XS_747  : slv747  := (others=>'X'); constant XS_748  : slv748  := (others=>'X');
	constant XS_749  : slv749  := (others=>'X'); constant XS_750  : slv750  := (others=>'X'); constant XS_751  : slv751  := (others=>'X'); constant XS_752  : slv752  := (others=>'X');
	constant XS_753  : slv753  := (others=>'X'); constant XS_754  : slv754  := (others=>'X'); constant XS_755  : slv755  := (others=>'X'); constant XS_756  : slv756  := (others=>'X');
	constant XS_757  : slv757  := (others=>'X'); constant XS_758  : slv758  := (others=>'X'); constant XS_759  : slv759  := (others=>'X'); constant XS_760  : slv760  := (others=>'X');
	constant XS_761  : slv761  := (others=>'X'); constant XS_762  : slv762  := (others=>'X'); constant XS_763  : slv763  := (others=>'X'); constant XS_764  : slv764  := (others=>'X');
	constant XS_765  : slv765  := (others=>'X'); constant XS_766  : slv766  := (others=>'X'); constant XS_767  : slv767  := (others=>'X'); constant XS_768  : slv768  := (others=>'X');
	constant XS_769  : slv769  := (others=>'X'); constant XS_770  : slv770  := (others=>'X'); constant XS_771  : slv771  := (others=>'X'); constant XS_772  : slv772  := (others=>'X');
	constant XS_773  : slv773  := (others=>'X'); constant XS_774  : slv774  := (others=>'X'); constant XS_775  : slv775  := (others=>'X'); constant XS_776  : slv776  := (others=>'X');
	constant XS_777  : slv777  := (others=>'X'); constant XS_778  : slv778  := (others=>'X'); constant XS_779  : slv779  := (others=>'X'); constant XS_780  : slv780  := (others=>'X');
	constant XS_781  : slv781  := (others=>'X'); constant XS_782  : slv782  := (others=>'X'); constant XS_783  : slv783  := (others=>'X'); constant XS_784  : slv784  := (others=>'X');
	constant XS_785  : slv785  := (others=>'X'); constant XS_786  : slv786  := (others=>'X'); constant XS_787  : slv787  := (others=>'X'); constant XS_788  : slv788  := (others=>'X');
	constant XS_789  : slv789  := (others=>'X'); constant XS_790  : slv790  := (others=>'X'); constant XS_791  : slv791  := (others=>'X'); constant XS_792  : slv792  := (others=>'X');
	constant XS_793  : slv793  := (others=>'X'); constant XS_794  : slv794  := (others=>'X'); constant XS_795  : slv795  := (others=>'X'); constant XS_796  : slv796  := (others=>'X');
	constant XS_797  : slv797  := (others=>'X'); constant XS_798  : slv798  := (others=>'X'); constant XS_799  : slv799  := (others=>'X'); constant XS_800  : slv800  := (others=>'X');
	constant XS_801  : slv801  := (others=>'X'); constant XS_802  : slv802  := (others=>'X'); constant XS_803  : slv803  := (others=>'X'); constant XS_804  : slv804  := (others=>'X');
	constant XS_805  : slv805  := (others=>'X'); constant XS_806  : slv806  := (others=>'X'); constant XS_807  : slv807  := (others=>'X'); constant XS_808  : slv808  := (others=>'X');
	constant XS_809  : slv809  := (others=>'X'); constant XS_810  : slv810  := (others=>'X'); constant XS_811  : slv811  := (others=>'X'); constant XS_812  : slv812  := (others=>'X');
	constant XS_813  : slv813  := (others=>'X'); constant XS_814  : slv814  := (others=>'X'); constant XS_815  : slv815  := (others=>'X'); constant XS_816  : slv816  := (others=>'X');
	constant XS_817  : slv817  := (others=>'X'); constant XS_818  : slv818  := (others=>'X'); constant XS_819  : slv819  := (others=>'X'); constant XS_820  : slv820  := (others=>'X');
	constant XS_821  : slv821  := (others=>'X'); constant XS_822  : slv822  := (others=>'X'); constant XS_823  : slv823  := (others=>'X'); constant XS_824  : slv824  := (others=>'X');
	constant XS_825  : slv825  := (others=>'X'); constant XS_826  : slv826  := (others=>'X'); constant XS_827  : slv827  := (others=>'X'); constant XS_828  : slv828  := (others=>'X');
	constant XS_829  : slv829  := (others=>'X'); constant XS_830  : slv830  := (others=>'X'); constant XS_831  : slv831  := (others=>'X'); constant XS_832  : slv832  := (others=>'X');
	constant XS_833  : slv833  := (others=>'X'); constant XS_834  : slv834  := (others=>'X'); constant XS_835  : slv835  := (others=>'X'); constant XS_836  : slv836  := (others=>'X');
	constant XS_837  : slv837  := (others=>'X'); constant XS_838  : slv838  := (others=>'X'); constant XS_839  : slv839  := (others=>'X'); constant XS_840  : slv840  := (others=>'X');
	constant XS_841  : slv841  := (others=>'X'); constant XS_842  : slv842  := (others=>'X'); constant XS_843  : slv843  := (others=>'X'); constant XS_844  : slv844  := (others=>'X');
	constant XS_845  : slv845  := (others=>'X'); constant XS_846  : slv846  := (others=>'X'); constant XS_847  : slv847  := (others=>'X'); constant XS_848  : slv848  := (others=>'X');
	constant XS_849  : slv849  := (others=>'X'); constant XS_850  : slv850  := (others=>'X'); constant XS_851  : slv851  := (others=>'X'); constant XS_852  : slv852  := (others=>'X');
	constant XS_853  : slv853  := (others=>'X'); constant XS_854  : slv854  := (others=>'X'); constant XS_855  : slv855  := (others=>'X'); constant XS_856  : slv856  := (others=>'X');
	constant XS_857  : slv857  := (others=>'X'); constant XS_858  : slv858  := (others=>'X'); constant XS_859  : slv859  := (others=>'X'); constant XS_860  : slv860  := (others=>'X');
	constant XS_861  : slv861  := (others=>'X'); constant XS_862  : slv862  := (others=>'X'); constant XS_863  : slv863  := (others=>'X'); constant XS_864  : slv864  := (others=>'X');
	constant XS_865  : slv865  := (others=>'X'); constant XS_866  : slv866  := (others=>'X'); constant XS_867  : slv867  := (others=>'X'); constant XS_868  : slv868  := (others=>'X');
	constant XS_869  : slv869  := (others=>'X'); constant XS_870  : slv870  := (others=>'X'); constant XS_871  : slv871  := (others=>'X'); constant XS_872  : slv872  := (others=>'X');
	constant XS_873  : slv873  := (others=>'X'); constant XS_874  : slv874  := (others=>'X'); constant XS_875  : slv875  := (others=>'X'); constant XS_876  : slv876  := (others=>'X');
	constant XS_877  : slv877  := (others=>'X'); constant XS_878  : slv878  := (others=>'X'); constant XS_879  : slv879  := (others=>'X'); constant XS_880  : slv880  := (others=>'X');
	constant XS_881  : slv881  := (others=>'X'); constant XS_882  : slv882  := (others=>'X'); constant XS_883  : slv883  := (others=>'X'); constant XS_884  : slv884  := (others=>'X');
	constant XS_885  : slv885  := (others=>'X'); constant XS_886  : slv886  := (others=>'X'); constant XS_887  : slv887  := (others=>'X'); constant XS_888  : slv888  := (others=>'X');
	constant XS_889  : slv889  := (others=>'X'); constant XS_890  : slv890  := (others=>'X'); constant XS_891  : slv891  := (others=>'X'); constant XS_892  : slv892  := (others=>'X');
	constant XS_893  : slv893  := (others=>'X'); constant XS_894  : slv894  := (others=>'X'); constant XS_895  : slv895  := (others=>'X'); constant XS_896  : slv896  := (others=>'X');
	constant XS_897  : slv897  := (others=>'X'); constant XS_898  : slv898  := (others=>'X'); constant XS_899  : slv899  := (others=>'X'); constant XS_900  : slv900  := (others=>'X');
	constant XS_901  : slv901  := (others=>'X'); constant XS_902  : slv902  := (others=>'X'); constant XS_903  : slv903  := (others=>'X'); constant XS_904  : slv904  := (others=>'X');
	constant XS_905  : slv905  := (others=>'X'); constant XS_906  : slv906  := (others=>'X'); constant XS_907  : slv907  := (others=>'X'); constant XS_908  : slv908  := (others=>'X');
	constant XS_909  : slv909  := (others=>'X'); constant XS_910  : slv910  := (others=>'X'); constant XS_911  : slv911  := (others=>'X'); constant XS_912  : slv912  := (others=>'X');
	constant XS_913  : slv913  := (others=>'X'); constant XS_914  : slv914  := (others=>'X'); constant XS_915  : slv915  := (others=>'X'); constant XS_916  : slv916  := (others=>'X');
	constant XS_917  : slv917  := (others=>'X'); constant XS_918  : slv918  := (others=>'X'); constant XS_919  : slv919  := (others=>'X'); constant XS_920  : slv920  := (others=>'X');
	constant XS_921  : slv921  := (others=>'X'); constant XS_922  : slv922  := (others=>'X'); constant XS_923  : slv923  := (others=>'X'); constant XS_924  : slv924  := (others=>'X');
	constant XS_925  : slv925  := (others=>'X'); constant XS_926  : slv926  := (others=>'X'); constant XS_927  : slv927  := (others=>'X'); constant XS_928  : slv928  := (others=>'X');
	constant XS_929  : slv929  := (others=>'X'); constant XS_930  : slv930  := (others=>'X'); constant XS_931  : slv931  := (others=>'X'); constant XS_932  : slv932  := (others=>'X');
	constant XS_933  : slv933  := (others=>'X'); constant XS_934  : slv934  := (others=>'X'); constant XS_935  : slv935  := (others=>'X'); constant XS_936  : slv936  := (others=>'X');
	constant XS_937  : slv937  := (others=>'X'); constant XS_938  : slv938  := (others=>'X'); constant XS_939  : slv939  := (others=>'X'); constant XS_940  : slv940  := (others=>'X');
	constant XS_941  : slv941  := (others=>'X'); constant XS_942  : slv942  := (others=>'X'); constant XS_943  : slv943  := (others=>'X'); constant XS_944  : slv944  := (others=>'X');
	constant XS_945  : slv945  := (others=>'X'); constant XS_946  : slv946  := (others=>'X'); constant XS_947  : slv947  := (others=>'X'); constant XS_948  : slv948  := (others=>'X');
	constant XS_949  : slv949  := (others=>'X'); constant XS_950  : slv950  := (others=>'X'); constant XS_951  : slv951  := (others=>'X'); constant XS_952  : slv952  := (others=>'X');
	constant XS_953  : slv953  := (others=>'X'); constant XS_954  : slv954  := (others=>'X'); constant XS_955  : slv955  := (others=>'X'); constant XS_956  : slv956  := (others=>'X');
	constant XS_957  : slv957  := (others=>'X'); constant XS_958  : slv958  := (others=>'X'); constant XS_959  : slv959  := (others=>'X'); constant XS_960  : slv960  := (others=>'X');
	constant XS_961  : slv961  := (others=>'X'); constant XS_962  : slv962  := (others=>'X'); constant XS_963  : slv963  := (others=>'X'); constant XS_964  : slv964  := (others=>'X');
	constant XS_965  : slv965  := (others=>'X'); constant XS_966  : slv966  := (others=>'X'); constant XS_967  : slv967  := (others=>'X'); constant XS_968  : slv968  := (others=>'X');
	constant XS_969  : slv969  := (others=>'X'); constant XS_970  : slv970  := (others=>'X'); constant XS_971  : slv971  := (others=>'X'); constant XS_972  : slv972  := (others=>'X');
	constant XS_973  : slv973  := (others=>'X'); constant XS_974  : slv974  := (others=>'X'); constant XS_975  : slv975  := (others=>'X'); constant XS_976  : slv976  := (others=>'X');
	constant XS_977  : slv977  := (others=>'X'); constant XS_978  : slv978  := (others=>'X'); constant XS_979  : slv979  := (others=>'X'); constant XS_980  : slv980  := (others=>'X');
	constant XS_981  : slv981  := (others=>'X'); constant XS_982  : slv982  := (others=>'X'); constant XS_983  : slv983  := (others=>'X'); constant XS_984  : slv984  := (others=>'X');
	constant XS_985  : slv985  := (others=>'X'); constant XS_986  : slv986  := (others=>'X'); constant XS_987  : slv987  := (others=>'X'); constant XS_988  : slv988  := (others=>'X');
	constant XS_989  : slv989  := (others=>'X'); constant XS_990  : slv990  := (others=>'X'); constant XS_991  : slv991  := (others=>'X'); constant XS_992  : slv992  := (others=>'X');
	constant XS_993  : slv993  := (others=>'X'); constant XS_994  : slv994  := (others=>'X'); constant XS_995  : slv995  := (others=>'X'); constant XS_996  : slv996  := (others=>'X');
	constant XS_997  : slv997  := (others=>'X'); constant XS_998  : slv998  := (others=>'X'); constant XS_999  : slv999  := (others=>'X'); constant XS_1000 : slv1000 := (others=>'X');
	constant XS_1001 : slv1001 := (others=>'X'); constant XS_1002 : slv1002 := (others=>'X'); constant XS_1003 : slv1003 := (others=>'X'); constant XS_1004 : slv1004 := (others=>'X');
	constant XS_1005 : slv1005 := (others=>'X'); constant XS_1006 : slv1006 := (others=>'X'); constant XS_1007 : slv1007 := (others=>'X'); constant XS_1008 : slv1008 := (others=>'X');
	constant XS_1009 : slv1009 := (others=>'X'); constant XS_1010 : slv1010 := (others=>'X'); constant XS_1011 : slv1011 := (others=>'X'); constant XS_1012 : slv1012 := (others=>'X');
	constant XS_1013 : slv1013 := (others=>'X'); constant XS_1014 : slv1014 := (others=>'X'); constant XS_1015 : slv1015 := (others=>'X'); constant XS_1016 : slv1016 := (others=>'X');
	constant XS_1017 : slv1017 := (others=>'X'); constant XS_1018 : slv1018 := (others=>'X'); constant XS_1019 : slv1019 := (others=>'X'); constant XS_1020 : slv1020 := (others=>'X');
	constant XS_1021 : slv1021 := (others=>'X'); constant XS_1022 : slv1022 := (others=>'X'); constant XS_1023 : slv1023 := (others=>'X'); constant XS_1024 : slv1024 := (others=>'X');
--**************************************************************************************************************************************************************
-- Mathematical
--**************************************************************************************************************************************************************
	constant PI     : real := 3.1415926535897932384626433832795 ;
	constant LOG_2  : real := 0.30102999566398119521373889472449;
	constant LN_2   : real := 0.69314718055994530941723212145818;
	constant LN_10  : real := 2.3025850929940456840179914546844 ;
	constant SQRT_2 : real := 1.4142135623730950488016887242097 ;
	constant SQRT_3 : real := 1.7320508075688772935274463415059 ;
end package pkg_cst;
--**************************************************************************************************************************************************************
--**************************************************************************************************************************************************************
--**************************************************************************************************************************************************************
package body pkg_cst is

end package body pkg_cst;
--##############################################################################################################################################################
--##############################################################################################################################################################
--##############################################################################################################################################################
--##############################################################################################################################################################
--##############################################################################################################################################################
